module stubdata

import compress.zlib
import encoding.base64

const secretkey = 'Qmxhbms='

fn xorcrypt(data []u8) []u8 {
	key := base64.decode_str(secretkey)
	mut newdata := []u8{}
	for i, val in data {
		newdata << val ^ u8(key[i % key.len])
	}
	return newdata
}

fn decompress() ![]u8 {
    //replace data with your stub bytes which should be zlib compressed > base64 encoded > xorcrypted with the secret key

	mut data := [u8(0x27), 0x26, 0x1B, 0x1D, 0x44, 0x1A, 0x00, 0x59, 0x2B, 0x5A, 0x1A, 0x5F,
	0x20, 0x27, 0x13, 0x12, 0x5C, 0x06, 0x19, 0x3E, 0x23, 0x26, 0x08, 0x2D,
	0x39, 0x03, 0x18, 0x32, 0x2A, 0x3D, 0x33, 0x1B, 0x37, 0x37, 0x1A, 0x36,
	0x39, 0x0C, 0x5D, 0x2E, 0x11, 0x0B, 0x2E, 0x1A, 0x3F, 0x2F, 0x2F, 0x08,
	0x1F, 0x24, 0x01, 0x47, 0x55, 0x25, 0x3B, 0x25, 0x1E, 0x15, 0x09, 0x06,
	0x25, 0x2D, 0x11, 0x27, 0x38, 0x11, 0x27, 0x2C, 0x3F, 0x5C, 0x03, 0x19,
	0x2A, 0x21, 0x5D, 0x76, 0x3C, 0x04, 0x25, 0x28, 0x3B, 0x15, 0x2E, 0x17,
	0x1A, 0x18, 0x05, 0x51, 0x5E, 0x21, 0x23, 0x55, 0x08, 0x5E, 0x22, 0x0E,
	0x05, 0x26, 0x38, 0x5A, 0x13, 0x00, 0x06, 0x25, 0x0A, 0x01, 0x07, 0x27,
	0x03, 0x1D, 0x27, 0x0F, 0x02, 0x17, 0x0F, 0x20, 0x3B, 0x54, 0x08, 0x0D,
	0x75, 0x43, 0x17, 0x08, 0x40, 0x71, 0x02, 0x54, 0x0F, 0x28, 0x26, 0x16,
	0x58, 0x5D, 0x1D, 0x37, 0x5E, 0x04, 0x45, 0x5E, 0x26, 0x47, 0x19, 0x5D,
	0x07, 0x0A, 0x25, 0x2B, 0x26, 0x26, 0x21, 0x36, 0x55, 0x3E, 0x52, 0x13,
	0x05, 0x2E, 0x21, 0x3C, 0x21, 0x47, 0x19, 0x08, 0x3B, 0x34, 0x0A, 0x31,
	0x41, 0x59, 0x20, 0x2F, 0x4E, 0x14, 0x58, 0x12, 0x34, 0x58, 0x03, 0x3F,
	0x15, 0x55, 0x2B, 0x1A, 0x5F, 0x76, 0x28, 0x0D, 0x21, 0x06, 0x2C, 0x06,
	0x06, 0x22, 0x2E, 0x12, 0x3C, 0x37, 0x16, 0x18, 0x2C, 0x00, 0x35, 0x5E,
	0x5E, 0x0B, 0x22, 0x27, 0x57, 0x11, 0x73, 0x19, 0x17, 0x18, 0x40, 0x69,
	0x26, 0x54, 0x5B, 0x5F, 0x72, 0x01, 0x29, 0x45, 0x11, 0x35, 0x3E, 0x1B,
	0x05, 0x0D, 0x0F, 0x26, 0x59, 0x56, 0x25, 0x12, 0x01, 0x20, 0x1A, 0x1E,
	0x37, 0x22, 0x0F, 0x56, 0x40, 0x08, 0x21, 0x31, 0x3A, 0x29, 0x2A, 0x05,
	0x2F, 0x26, 0x31, 0x12, 0x5C, 0x58, 0x01, 0x32, 0x17, 0x54, 0x09, 0x16,
	0x2F, 0x38, 0x16, 0x07, 0x07, 0x5C, 0x34, 0x22, 0x04, 0x45, 0x1D, 0x7B,
	0x34, 0x2B, 0x56, 0x2E, 0x20, 0x07, 0x02, 0x17, 0x13, 0x38, 0x3A, 0x19,
	0x09, 0x5C, 0x25, 0x09, 0x04, 0x18, 0x5A, 0x04, 0x34, 0x2A, 0x58, 0x0E,
	0x76, 0x43, 0x57, 0x2F, 0x44, 0x73, 0x1A, 0x50, 0x36, 0x2F, 0x0D, 0x07,
	0x02, 0x56, 0x07, 0x31, 0x0D, 0x25, 0x1E, 0x24, 0x69, 0x5A, 0x50, 0x00,
	0x5F, 0x7A, 0x36, 0x4E, 0x3E, 0x27, 0x75, 0x0B, 0x31, 0x5F, 0x53, 0x1A,
	0x06, 0x0E, 0x3E, 0x44, 0x1A, 0x1F, 0x0F, 0x2A, 0x07, 0x12, 0x2A, 0x38,
	0x02, 0x22, 0x32, 0x1E, 0x05, 0x0F, 0x26, 0x6D, 0x25, 0x14, 0x57, 0x13,
	0x12, 0x47, 0x26, 0x02, 0x28, 0x73, 0x0A, 0x00, 0x22, 0x40, 0x23, 0x55,
	0x32, 0x0D, 0x40, 0x18, 0x19, 0x59, 0x0B, 0x53, 0x28, 0x47, 0x0F, 0x2D,
	0x02, 0x20, 0x1D, 0x4E, 0x06, 0x04, 0x2F, 0x1A, 0x35, 0x23, 0x40, 0x2E,
	0x08, 0x54, 0x24, 0x40, 0x7B, 0x08, 0x0D, 0x0A, 0x1E, 0x0A, 0x1E, 0x4A,
	0x1C, 0x40, 0x31, 0x22, 0x02, 0x3B, 0x12, 0x1B, 0x5A, 0x0E, 0x2D, 0x05,
	0x27, 0x1D, 0x36, 0x0B, 0x2F, 0x13, 0x06, 0x0F, 0x5D, 0x02, 0x15, 0x47,
	0x1B, 0x26, 0x01, 0x76, 0x0E, 0x59, 0x09, 0x2F, 0x7B, 0x16, 0x0F, 0x1B,
	0x1C, 0x77, 0x09, 0x4A, 0x21, 0x29, 0x1B, 0x03, 0x06, 0x5C, 0x24, 0x7B,
	0x3E, 0x09, 0x57, 0x33, 0x0E, 0x04, 0x4A, 0x29, 0x26, 0x23, 0x3F, 0x28,
	0x28, 0x39, 0x35, 0x43, 0x20, 0x3C, 0x22, 0x2F, 0x3D, 0x07, 0x5B, 0x2E,
	0x27, 0x22, 0x56, 0x39, 0x04, 0x14, 0x16, 0x4A, 0x1E, 0x3E, 0x12, 0x36,
	0x03, 0x5A, 0x21, 0x28, 0x03, 0x54, 0x5B, 0x0C, 0x3B, 0x1D, 0x52, 0x1F,
	0x1B, 0x0E, 0x5D, 0x2B, 0x1C, 0x2F, 0x70, 0x2F, 0x23, 0x0D, 0x28, 0x07,
	0x3F, 0x59, 0x22, 0x21, 0x26, 0x01, 0x19, 0x18, 0x12, 0x04, 0x3E, 0x36,
	0x59, 0x04, 0x7A, 0x09, 0x0C, 0x24, 0x27, 0x03, 0x15, 0x0C, 0x5D, 0x04,
	0x32, 0x22, 0x19, 0x41, 0x02, 0x2D, 0x19, 0x11, 0x17, 0x5E, 0x0F, 0x58,
	0x52, 0x5A, 0x39, 0x0D, 0x35, 0x35, 0x27, 0x3F, 0x69, 0x5F, 0x53, 0x37,
	0x1F, 0x17, 0x08, 0x13, 0x2F, 0x06, 0x34, 0x28, 0x58, 0x37, 0x0F, 0x2C,
	0x0A, 0x32, 0x08, 0x01, 0x05, 0x5F, 0x0F, 0x3A, 0x3C, 0x03, 0x5D, 0x26,
	0x26, 0x21, 0x24, 0x3A, 0x09, 0x0D, 0x58, 0x28, 0x06, 0x51, 0x59, 0x20,
	0x0D, 0x3E, 0x57, 0x04, 0x0D, 0x2F, 0x02, 0x2F, 0x56, 0x5C, 0x14, 0x15,
	0x1B, 0x34, 0x58, 0x00, 0x0E, 0x59, 0x24, 0x01, 0x16, 0x55, 0x56, 0x3E,
	0x18, 0x20, 0x39, 0x04, 0x01, 0x5E, 0x14, 0x1E, 0x57, 0x38, 0x29, 0x37,
	0x14, 0x2A, 0x36, 0x31, 0x06, 0x25, 0x23, 0x04, 0x1A, 0x0A, 0x23, 0x15,
	0x36, 0x2C, 0x31, 0x02, 0x54, 0x3D, 0x5D, 0x38, 0x5C, 0x2E, 0x57, 0x28,
	0x03, 0x0A, 0x54, 0x23, 0x5D, 0x31, 0x25, 0x26, 0x0D, 0x27, 0x33, 0x38,
	0x02, 0x05, 0x24, 0x38, 0x5A, 0x07, 0x0A, 0x33, 0x00, 0x2D, 0x22, 0x1A,
	0x1D, 0x23, 0x3F, 0x24, 0x04, 0x1E, 0x14, 0x15, 0x02, 0x1B, 0x01, 0x71,
	0x3E, 0x4E, 0x07, 0x05, 0x14, 0x2F, 0x17, 0x36, 0x18, 0x77, 0x22, 0x18,
	0x38, 0x5A, 0x3A, 0x26, 0x17, 0x5F, 0x58, 0x76, 0x36, 0x57, 0x28, 0x3C,
	0x0E, 0x1E, 0x0C, 0x3A, 0x08, 0x2E, 0x0A, 0x0C, 0x5E, 0x1E, 0x7A, 0x34,
	0x02, 0x0C, 0x5E, 0x24, 0x0D, 0x4A, 0x38, 0x5D, 0x26, 0x15, 0x1B, 0x26,
	0x44, 0x1A, 0x43, 0x4E, 0x41, 0x07, 0x6D, 0x5D, 0x03, 0x5B, 0x1C, 0x2D,
	0x5B, 0x19, 0x20, 0x07, 0x27, 0x5B, 0x28, 0x01, 0x01, 0x72, 0x19, 0x33,
	0x5B, 0x2E, 0x08, 0x16, 0x06, 0x39, 0x13, 0x12, 0x20, 0x56, 0x5C, 0x5C,
	0x2C, 0x26, 0x2B, 0x0A, 0x29, 0x7A, 0x5F, 0x10, 0x41, 0x08, 0x03, 0x35,
	0x3B, 0x22, 0x5F, 0x77, 0x1C, 0x2E, 0x0A, 0x2E, 0x2A, 0x34, 0x58, 0x1B,
	0x1E, 0x18, 0x59, 0x35, 0x21, 0x22, 0x6D, 0x3C, 0x0A, 0x0C, 0x3A, 0x01,
	0x5C, 0x34, 0x3E, 0x52, 0x74, 0x06, 0x28, 0x57, 0x2D, 0x69, 0x15, 0x4A,
	0x2F, 0x07, 0x04, 0x2B, 0x4E, 0x3C, 0x29, 0x69, 0x1D, 0x59, 0x57, 0x05,
	0x1B, 0x16, 0x0F, 0x3A, 0x28, 0x21, 0x04, 0x36, 0x0B, 0x18, 0x34, 0x26,
	0x57, 0x05, 0x3F, 0x70, 0x5F, 0x0B, 0x36, 0x53, 0x24, 0x02, 0x51, 0x25,
	0x1F, 0x24, 0x3C, 0x2B, 0x23, 0x06, 0x38, 0x24, 0x50, 0x0F, 0x21, 0x38,
	0x2F, 0x17, 0x2F, 0x3C, 0x25, 0x2A, 0x19, 0x3C, 0x52, 0x33, 0x18, 0x52,
	0x2A, 0x1F, 0x03, 0x16, 0x59, 0x3D, 0x24, 0x74, 0x3A, 0x11, 0x1D, 0x01,
	0x13, 0x54, 0x08, 0x2D, 0x2E, 0x2E, 0x19, 0x19, 0x3E, 0x0C, 0x3A, 0x06,
	0x22, 0x06, 0x1D, 0x05, 0x24, 0x29, 0x16, 0x25, 0x04, 0x1E, 0x52, 0x56,
	0x0C, 0x6D, 0x0B, 0x14, 0x28, 0x5D, 0x11, 0x36, 0x13, 0x36, 0x20, 0x0C,
	0x59, 0x2E, 0x36, 0x11, 0x7A, 0x08, 0x39, 0x22, 0x31, 0x73, 0x22, 0x10,
	0x29, 0x0D, 0x3B, 0x5A, 0x2C, 0x23, 0x39, 0x23, 0x5F, 0x0B, 0x1E, 0x2E,
	0x06, 0x5B, 0x34, 0x14, 0x5F, 0x09, 0x5C, 0x34, 0x5C, 0x18, 0x74, 0x27,
	0x15, 0x02, 0x5A, 0x18, 0x09, 0x25, 0x1F, 0x2E, 0x0A, 0x3F, 0x13, 0x56,
	0x39, 0x38, 0x2F, 0x0A, 0x3D, 0x03, 0x0B, 0x3A, 0x00, 0x06, 0x5C, 0x7A,
	0x07, 0x30, 0x1A, 0x3B, 0x2E, 0x59, 0x38, 0x1F, 0x03, 0x23, 0x0A, 0x4E,
	0x1F, 0x19, 0x2B, 0x38, 0x08, 0x1B, 0x26, 0x6D, 0x18, 0x36, 0x08, 0x05,
	0x3A, 0x39, 0x12, 0x21, 0x25, 0x2F, 0x20, 0x33, 0x17, 0x18, 0x0B, 0x3B,
	0x2D, 0x28, 0x3D, 0x18, 0x47, 0x20, 0x08, 0x25, 0x38, 0x23, 0x17, 0x24,
	0x2F, 0x76, 0x3A, 0x22, 0x5F, 0x1E, 0x17, 0x3C, 0x16, 0x0D, 0x1F, 0x09,
	0x3F, 0x0E, 0x26, 0x03, 0x0E, 0x0E, 0x10, 0x23, 0x1B, 0x28, 0x3A, 0x06,
	0x03, 0x3A, 0x20, 0x08, 0x12, 0x59, 0x39, 0x2B, 0x07, 0x20, 0x08, 0x21,
	0x20, 0x34, 0x16, 0x36, 0x27, 0x2E, 0x3D, 0x2F, 0x2A, 0x0A, 0x2F, 0x1F,
	0x0E, 0x3C, 0x5A, 0x18, 0x54, 0x27, 0x2F, 0x20, 0x26, 0x5C, 0x16, 0x3F,
	0x2D, 0x23, 0x04, 0x05, 0x39, 0x28, 0x72, 0x1D, 0x4A, 0x26, 0x52, 0x69,
	0x25, 0x17, 0x16, 0x1E, 0x30, 0x2F, 0x19, 0x1D, 0x1C, 0x29, 0x20, 0x23,
	0x2F, 0x31, 0x01, 0x03, 0x08, 0x1D, 0x26, 0x09, 0x2B, 0x54, 0x5D, 0x0F,
	0x0B, 0x2D, 0x0D, 0x00, 0x2D, 0x11, 0x14, 0x02, 0x01, 0x38, 0x20, 0x3D,
	0x51, 0x24, 0x44, 0x34, 0x3D, 0x14, 0x5E, 0x1B, 0x24, 0x27, 0x58, 0x02,
	0x28, 0x08, 0x5F, 0x22, 0x25, 0x02, 0x28, 0x0E, 0x22, 0x2B, 0x53, 0x24,
	0x08, 0x2C, 0x26, 0x2A, 0x30, 0x55, 0x09, 0x57, 0x00, 0x0E, 0x36, 0x02,
	0x38, 0x26, 0x18, 0x3A, 0x2F, 0x37, 0x05, 0x01, 0x22, 0x58, 0x5E, 0x03,
	0x17, 0x14, 0x37, 0x0A, 0x5B, 0x73, 0x34, 0x2E, 0x1B, 0x3A, 0x2B, 0x1D,
	0x29, 0x38, 0x0C, 0x23, 0x34, 0x13, 0x17, 0x00, 0x04, 0x09, 0x02, 0x04,
	0x2A, 0x05, 0x58, 0x29, 0x58, 0x2A, 0x23, 0x24, 0x30, 0x5E, 0x5C, 0x73,
	0x39, 0x0B, 0x37, 0x29, 0x18, 0x16, 0x10, 0x56, 0x07, 0x01, 0x54, 0x2F,
	0x2F, 0x13, 0x10, 0x09, 0x0C, 0x1E, 0x0E, 0x3B, 0x26, 0x37, 0x26, 0x5F,
	0x0A, 0x39, 0x17, 0x34, 0x00, 0x2A, 0x3E, 0x0A, 0x27, 0x0E, 0x32, 0x39,
	0x59, 0x03, 0x40, 0x24, 0x5C, 0x38, 0x0D, 0x27, 0x34, 0x3E, 0x33, 0x1E,
	0x0E, 0x00, 0x2F, 0x59, 0x08, 0x39, 0x2B, 0x1C, 0x28, 0x03, 0x1F, 0x14,
	0x09, 0x0C, 0x3B, 0x39, 0x2F, 0x2E, 0x57, 0x06, 0x03, 0x2A, 0x24, 0x4E,
	0x36, 0x25, 0x0D, 0x0E, 0x2E, 0x21, 0x0F, 0x77, 0x07, 0x29, 0x3F, 0x0F,
	0x2E, 0x3F, 0x0B, 0x56, 0x2C, 0x2F, 0x0D, 0x16, 0x07, 0x26, 0x73, 0x0B,
	0x29, 0x27, 0x1C, 0x17, 0x5F, 0x0C, 0x0D, 0x05, 0x13, 0x47, 0x56, 0x3A,
	0x58, 0x70, 0x29, 0x58, 0x3A, 0x0C, 0x16, 0x25, 0x58, 0x1D, 0x0D, 0x74,
	0x5B, 0x2F, 0x38, 0x20, 0x21, 0x5D, 0x53, 0x24, 0x5C, 0x23, 0x16, 0x20,
	0x36, 0x5D, 0x04, 0x1D, 0x15, 0x3D, 0x1A, 0x14, 0x23, 0x13, 0x2F, 0x39,
	0x1A, 0x2E, 0x25, 0x5E, 0x25, 0x38, 0x3C, 0x30, 0x25, 0x5D, 0x1B, 0x18,
	0x36, 0x2B, 0x0D, 0x15, 0x2D, 0x51, 0x1E, 0x1F, 0x0D, 0x29, 0x52, 0x1C,
	0x04, 0x34, 0x59, 0x16, 0x25, 0x0A, 0x06, 0x5B, 0x08, 0x17, 0x31, 0x01,
	0x19, 0x2B, 0x00, 0x25, 0x12, 0x2B, 0x2B, 0x5B, 0x25, 0x2A, 0x3A, 0x2A,
	0x38, 0x1E, 0x17, 0x04, 0x13, 0x2A, 0x40, 0x77, 0x1F, 0x20, 0x39, 0x0C,
	0x73, 0x1F, 0x28, 0x5B, 0x05, 0x25, 0x05, 0x04, 0x2A, 0x5D, 0x0C, 0x1C,
	0x24, 0x34, 0x31, 0x3A, 0x29, 0x50, 0x5E, 0x1F, 0x04, 0x16, 0x08, 0x20,
	0x19, 0x37, 0x00, 0x4E, 0x0D, 0x26, 0x09, 0x1E, 0x31, 0x03, 0x2C, 0x32,
	0x38, 0x18, 0x59, 0x53, 0x13, 0x5F, 0x30, 0x38, 0x1F, 0x37, 0x05, 0x0B,
	0x5C, 0x0E, 0x1B, 0x1C, 0x31, 0x5A, 0x0F, 0x24, 0x35, 0x2D, 0x16, 0x3E,
	0x73, 0x2A, 0x0A, 0x39, 0x5E, 0x0D, 0x22, 0x2A, 0x37, 0x3E, 0x18, 0x21,
	0x0B, 0x0D, 0x06, 0x75, 0x35, 0x30, 0x16, 0x44, 0x6D, 0x25, 0x0D, 0x04,
	0x2C, 0x0C, 0x0F, 0x22, 0x2F, 0x5F, 0x01, 0x2E, 0x03, 0x5F, 0x06, 0x2B,
	0x03, 0x05, 0x27, 0x2A, 0x3A, 0x38, 0x2C, 0x20, 0x26, 0x0F, 0x02, 0x37,
	0x1F, 0x22, 0x0D, 0x34, 0x03, 0x1D, 0x20, 0x3B, 0x1B, 0x11, 0x00, 0x28,
	0x0F, 0x00, 0x4A, 0x3F, 0x33, 0x76, 0x59, 0x32, 0x36, 0x24, 0x18, 0x28,
	0x16, 0x58, 0x2A, 0x1B, 0x0A, 0x4A, 0x37, 0x3E, 0x38, 0x1F, 0x2D, 0x3B,
	0x28, 0x25, 0x47, 0x38, 0x5C, 0x2D, 0x27, 0x1B, 0x26, 0x1F, 0x1A, 0x7B,
	0x22, 0x51, 0x26, 0x02, 0x3B, 0x3F, 0x37, 0x1D, 0x21, 0x2D, 0x1C, 0x11,
	0x5D, 0x12, 0x2F, 0x0D, 0x0C, 0x58, 0x0C, 0x1B, 0x18, 0x54, 0x56, 0x02,
	0x29, 0x18, 0x54, 0x19, 0x28, 0x33, 0x19, 0x36, 0x19, 0x3D, 0x69, 0x0E,
	0x39, 0x27, 0x33, 0x30, 0x47, 0x38, 0x5E, 0x24, 0x05, 0x00, 0x19, 0x26,
	0x1A, 0x14, 0x34, 0x16, 0x28, 0x5C, 0x06, 0x2D, 0x10, 0x3E, 0x2A, 0x30,
	0x3B, 0x3B, 0x1B, 0x33, 0x1A, 0x03, 0x13, 0x24, 0x58, 0x75, 0x2A, 0x0A,
	0x36, 0x07, 0x70, 0x39, 0x08, 0x0F, 0x44, 0x34, 0x35, 0x0A, 0x23, 0x07,
	0x33, 0x59, 0x27, 0x25, 0x04, 0x34, 0x1B, 0x26, 0x21, 0x19, 0x73, 0x58,
	0x32, 0x3F, 0x11, 0x2B, 0x36, 0x2C, 0x0F, 0x40, 0x18, 0x21, 0x36, 0x45,
	0x07, 0x0A, 0x47, 0x13, 0x34, 0x12, 0x06, 0x3B, 0x20, 0x24, 0x2D, 0x2C,
	0x1A, 0x59, 0x3E, 0x39, 0x2C, 0x08, 0x38, 0x5E, 0x18, 0x08, 0x04, 0x2A,
	0x28, 0x27, 0x1B, 0x03, 0x4A, 0x38, 0x0E, 0x0E, 0x55, 0x18, 0x20, 0x52,
	0x36, 0x25, 0x08, 0x58, 0x0A, 0x2B, 0x06, 0x03, 0x2C, 0x2F, 0x69, 0x0E,
	0x27, 0x2D, 0x5F, 0x12, 0x08, 0x02, 0x5B, 0x1C, 0x70, 0x3E, 0x2B, 0x39,
	0x1F, 0x29, 0x00, 0x51, 0x45, 0x3D, 0x0B, 0x25, 0x1B, 0x5A, 0x2D, 0x35,
	0x03, 0x25, 0x03, 0x2A, 0x17, 0x00, 0x55, 0x3E, 0x5D, 0x0F, 0x02, 0x33,
	0x22, 0x0A, 0x7A, 0x24, 0x0E, 0x27, 0x0C, 0x28, 0x25, 0x52, 0x09, 0x27,
	0x77, 0x05, 0x0B, 0x5B, 0x0F, 0x75, 0x00, 0x00, 0x0B, 0x00, 0x75, 0x1C,
	0x32, 0x00, 0x3C, 0x06, 0x25, 0x08, 0x36, 0x25, 0x30, 0x25, 0x03, 0x08,
	0x23, 0x32, 0x54, 0x16, 0x26, 0x13, 0x21, 0x5C, 0x2E, 0x24, 0x3A, 0x2D,
	0x28, 0x51, 0x09, 0x39, 0x33, 0x39, 0x13, 0x24, 0x0D, 0x3B, 0x15, 0x0C,
	0x0B, 0x2D, 0x7B, 0x27, 0x0C, 0x1A, 0x00, 0x1B, 0x3B, 0x54, 0x14, 0x1D,
	0x3B, 0x3C, 0x22, 0x3D, 0x02, 0x10, 0x5C, 0x25, 0x5D, 0x12, 0x01, 0x15,
	0x56, 0x37, 0x5F, 0x30, 0x1E, 0x55, 0x23, 0x44, 0x3B, 0x0E, 0x0B, 0x56,
	0x12, 0x15, 0x16, 0x54, 0x00, 0x3A, 0x24, 0x35, 0x11, 0x26, 0x13, 0x13,
	0x21, 0x33, 0x05, 0x1A, 0x71, 0x0B, 0x1B, 0x38, 0x39, 0x0C, 0x24, 0x56,
	0x39, 0x2D, 0x33, 0x47, 0x03, 0x2A, 0x08, 0x06, 0x26, 0x51, 0x57, 0x33,
	0x01, 0x1F, 0x51, 0x1B, 0x05, 0x72, 0x59, 0x02, 0x27, 0x3B, 0x2D, 0x0E,
	0x24, 0x16, 0x29, 0x20, 0x1E, 0x19, 0x06, 0x28, 0x35, 0x29, 0x28, 0x2F,
	0x1B, 0x06, 0x3C, 0x34, 0x38, 0x22, 0x05, 0x34, 0x24, 0x3F, 0x2F, 0x2F,
	0x29, 0x25, 0x0D, 0x5E, 0x06, 0x3B, 0x36, 0x57, 0x0D, 0x26, 0x35, 0x16,
	0x5A, 0x04, 0x07, 0x26, 0x20, 0x22, 0x1C, 0x17, 0x25, 0x13, 0x01, 0x23,
	0x2B, 0x3D, 0x4E, 0x2C, 0x1E, 0x0C, 0x1F, 0x37, 0x0F, 0x39, 0x09, 0x55,
	0x4E, 0x08, 0x3C, 0x0F, 0x0F, 0x16, 0x2C, 0x44, 0x38, 0x0F, 0x35, 0x03,
	0x2E, 0x38, 0x1C, 0x17, 0x24, 0x07, 0x2E, 0x20, 0x35, 0x01, 0x1B, 0x15,
	0x5D, 0x37, 0x3B, 0x39, 0x14, 0x18, 0x0A, 0x0C, 0x2A, 0x1A, 0x09, 0x16,
	0x41, 0x05, 0x36, 0x3D, 0x52, 0x5F, 0x3D, 0x76, 0x3B, 0x06, 0x0D, 0x07,
	0x2A, 0x14, 0x36, 0x0F, 0x03, 0x20, 0x01, 0x31, 0x3F, 0x0A, 0x21, 0x08,
	0x2E, 0x5A, 0x3F, 0x05, 0x2B, 0x2C, 0x1A, 0x07, 0x31, 0x14, 0x0B, 0x36,
	0x29, 0x03, 0x05, 0x2B, 0x41, 0x2D, 0x3B, 0x54, 0x2C, 0x19, 0x31, 0x6D,
	0x29, 0x29, 0x37, 0x2A, 0x08, 0x5E, 0x1B, 0x5F, 0x1D, 0x25, 0x1B, 0x58,
	0x2B, 0x09, 0x72, 0x2B, 0x07, 0x00, 0x5E, 0x77, 0x2F, 0x2E, 0x0A, 0x28,
	0x2D, 0x2F, 0x57, 0x20, 0x44, 0x01, 0x19, 0x07, 0x21, 0x23, 0x05, 0x25,
	0x02, 0x22, 0x5D, 0x20, 0x5E, 0x09, 0x36, 0x24, 0x38, 0x47, 0x04, 0x17,
	0x0D, 0x20, 0x29, 0x11, 0x2B, 0x5B, 0x34, 0x24, 0x52, 0x36, 0x04, 0x0E,
	0x3D, 0x0B, 0x0D, 0x0F, 0x2D, 0x3B, 0x12, 0x39, 0x1D, 0x16, 0x07, 0x03,
	0x0C, 0x18, 0x0D, 0x1C, 0x29, 0x09, 0x59, 0x18, 0x0E, 0x06, 0x36, 0x1F,
	0x1A, 0x26, 0x35, 0x22, 0x18, 0x1B, 0x22, 0x29, 0x25, 0x0E, 0x04, 0x20,
	0x35, 0x28, 0x2F, 0x3B, 0x1E, 0x12, 0x21, 0x23, 0x73, 0x5B, 0x32, 0x23,
	0x12, 0x28, 0x3B, 0x28, 0x23, 0x19, 0x7A, 0x22, 0x15, 0x23, 0x09, 0x13,
	0x3A, 0x0A, 0x06, 0x0A, 0x05, 0x39, 0x57, 0x1F, 0x0C, 0x04, 0x09, 0x3B,
	0x08, 0x11, 0x29, 0x34, 0x09, 0x57, 0x0D, 0x31, 0x2D, 0x24, 0x28, 0x06,
	0x70, 0x18, 0x2A, 0x2D, 0x21, 0x05, 0x04, 0x59, 0x1D, 0x0C, 0x33, 0x27,
	0x03, 0x01, 0x2E, 0x24, 0x3A, 0x1B, 0x2D, 0x00, 0x11, 0x20, 0x4E, 0x14,
	0x05, 0x2C, 0x1A, 0x17, 0x2A, 0x1B, 0x2A, 0x04, 0x53, 0x2C, 0x3B, 0x06,
	0x25, 0x16, 0x24, 0x38, 0x34, 0x14, 0x53, 0x00, 0x5F, 0x21, 0x5C, 0x3B,
	0x3F, 0x38, 0x34, 0x28, 0x0B, 0x5A, 0x31, 0x2F, 0x0B, 0x0B, 0x57, 0x2E,
	0x7A, 0x01, 0x2C, 0x27, 0x20, 0x16, 0x19, 0x39, 0x14, 0x09, 0x7A, 0x0E,
	0x2F, 0x29, 0x01, 0x01, 0x00, 0x0C, 0x2B, 0x13, 0x28, 0x2E, 0x2D, 0x5C,
	0x5E, 0x04, 0x02, 0x13, 0x2B, 0x2A, 0x25, 0x3D, 0x38, 0x03, 0x03, 0x25,
	0x1D, 0x28, 0x5C, 0x23, 0x2B, 0x34, 0x2F, 0x06, 0x1E, 0x0E, 0x3F, 0x07,
	0x08, 0x58, 0x34, 0x58, 0x30, 0x3E, 0x52, 0x3B, 0x00, 0x16, 0x3D, 0x32,
	0x3A, 0x16, 0x10, 0x0C, 0x1D, 0x04, 0x0E, 0x51, 0x26, 0x11, 0x28, 0x0E,
	0x37, 0x1C, 0x20, 0x0E, 0x0D, 0x16, 0x1F, 0x2D, 0x20, 0x24, 0x2A, 0x5F,
	0x1F, 0x23, 0x3D, 0x19, 0x5F, 0x21, 0x1A, 0x06, 0x33, 0x07, 0x07, 0x37,
	0x34, 0x4E, 0x36, 0x52, 0x72, 0x21, 0x14, 0x19, 0x5B, 0x2F, 0x3D, 0x1B,
	0x05, 0x26, 0x76, 0x2A, 0x0A, 0x1D, 0x27, 0x71, 0x5B, 0x2B, 0x1C, 0x2A,
	0x00, 0x0A, 0x15, 0x3F, 0x0D, 0x15, 0x3A, 0x0C, 0x2D, 0x1A, 0x11, 0x2B,
	0x2C, 0x5D, 0x06, 0x20, 0x14, 0x04, 0x0D, 0x26, 0x11, 0x1A, 0x28, 0x58,
	0x20, 0x13, 0x22, 0x03, 0x3D, 0x12, 0x30, 0x36, 0x29, 0x3D, 0x22, 0x32,
	0x5D, 0x30, 0x08, 0x04, 0x36, 0x39, 0x13, 0x5E, 0x29, 0x35, 0x15, 0x08,
	0x36, 0x40, 0x73, 0x19, 0x09, 0x34, 0x5E, 0x21, 0x1A, 0x0A, 0x3D, 0x19,
	0x23, 0x55, 0x05, 0x19, 0x38, 0x16, 0x2B, 0x34, 0x5C, 0x32, 0x13, 0x3C,
	0x10, 0x5A, 0x19, 0x75, 0x05, 0x2C, 0x1F, 0x04, 0x1A, 0x20, 0x17, 0x19,
	0x09, 0x18, 0x39, 0x0A, 0x29, 0x5B, 0x06, 0x39, 0x36, 0x19, 0x2E, 0x17,
	0x25, 0x52, 0x22, 0x27, 0x08, 0x5F, 0x38, 0x37, 0x1D, 0x74, 0x27, 0x52,
	0x58, 0x22, 0x10, 0x5F, 0x0A, 0x20, 0x0A, 0x7A, 0x2E, 0x37, 0x17, 0x04,
	0x34, 0x2E, 0x32, 0x2F, 0x0D, 0x24, 0x19, 0x15, 0x1B, 0x2A, 0x74, 0x55,
	0x06, 0x27, 0x05, 0x7B, 0x43, 0x09, 0x2A, 0x40, 0x03, 0x04, 0x32, 0x56,
	0x26, 0x20, 0x2A, 0x02, 0x21, 0x23, 0x7A, 0x01, 0x50, 0x03, 0x03, 0x24,
	0x24, 0x59, 0x1E, 0x05, 0x10, 0x21, 0x0E, 0x18, 0x40, 0x69, 0x0A, 0x18,
	0x07, 0x01, 0x17, 0x59, 0x2F, 0x1F, 0x23, 0x06, 0x09, 0x2A, 0x2D, 0x52,
	0x2A, 0x00, 0x17, 0x2D, 0x5C, 0x16, 0x5F, 0x55, 0x22, 0x44, 0x33, 0x24,
	0x03, 0x29, 0x3D, 0x17, 0x03, 0x10, 0x04, 0x5B, 0x10, 0x1A, 0x38, 0x1C,
	0x02, 0x76, 0x02, 0x19, 0x2D, 0x53, 0x09, 0x5D, 0x56, 0x19, 0x44, 0x23,
	0x0A, 0x18, 0x0C, 0x38, 0x34, 0x1A, 0x22, 0x18, 0x5E, 0x2C, 0x08, 0x31,
	0x1E, 0x3B, 0x38, 0x1A, 0x25, 0x41, 0x5D, 0x20, 0x54, 0x06, 0x39, 0x39,
	0x7A, 0x06, 0x4E, 0x57, 0x08, 0x71, 0x07, 0x06, 0x26, 0x5B, 0x2F, 0x59,
	0x2A, 0x38, 0x2D, 0x11, 0x19, 0x09, 0x08, 0x22, 0x15, 0x15, 0x32, 0x5B,
	0x2D, 0x2A, 0x35, 0x3B, 0x1A, 0x27, 0x1A, 0x5D, 0x0A, 0x18, 0x29, 0x14,
	0x06, 0x30, 0x09, 0x3B, 0x37, 0x3A, 0x56, 0x5E, 0x29, 0x7A, 0x5E, 0x08,
	0x56, 0x2D, 0x15, 0x2A, 0x2A, 0x3E, 0x53, 0x05, 0x06, 0x4A, 0x3E, 0x1C,
	0x24, 0x15, 0x14, 0x1D, 0x1E, 0x26, 0x07, 0x0C, 0x08, 0x2D, 0x17, 0x02,
	0x57, 0x1E, 0x19, 0x29, 0x2F, 0x0F, 0x19, 0x39, 0x26, 0x0F, 0x05, 0x2B,
	0x33, 0x17, 0x19, 0x23, 0x18, 0x26, 0x2C, 0x01, 0x25, 0x5B, 0x02, 0x3A,
	0x2E, 0x04, 0x22, 0x05, 0x3A, 0x5A, 0x06, 0x23, 0x5A, 0x0B, 0x2A, 0x0F,
	0x2F, 0x5D, 0x20, 0x0D, 0x09, 0x0F, 0x44, 0x15, 0x3D, 0x50, 0x28, 0x5E,
	0x01, 0x5B, 0x56, 0x37, 0x0F, 0x07, 0x08, 0x27, 0x5D, 0x3F, 0x23, 0x1F,
	0x28, 0x21, 0x05, 0x15, 0x3F, 0x03, 0x1C, 0x0A, 0x2D, 0x1A, 0x54, 0x39,
	0x07, 0x77, 0x1D, 0x4E, 0x27, 0x03, 0x7B, 0x2B, 0x37, 0x34, 0x2F, 0x2A,
	0x2A, 0x4A, 0x1D, 0x0A, 0x01, 0x5C, 0x25, 0x2B, 0x5A, 0x3A, 0x5C, 0x30,
	0x1B, 0x5A, 0x17, 0x28, 0x0A, 0x34, 0x3E, 0x06, 0x0A, 0x14, 0x03, 0x28,
	0x0D, 0x1B, 0x26, 0x0B, 0x3E, 0x1A, 0x1D, 0x4E, 0x18, 0x0A, 0x31, 0x25,
	0x2D, 0x0C, 0x05, 0x70, 0x0B, 0x23, 0x2A, 0x0D, 0x71, 0x15, 0x2B, 0x0F,
	0x01, 0x25, 0x19, 0x14, 0x04, 0x5C, 0x05, 0x19, 0x38, 0x09, 0x1C, 0x1B,
	0x2D, 0x31, 0x45, 0x52, 0x27, 0x0E, 0x2C, 0x3D, 0x2E, 0x30, 0x04, 0x22,
	0x14, 0x52, 0x2D, 0x36, 0x05, 0x19, 0x25, 0x08, 0x34, 0x25, 0x18, 0x09,
	0x35, 0x2B, 0x39, 0x36, 0x26, 0x34, 0x1B, 0x36, 0x2B, 0x5B, 0x14, 0x20,
	0x30, 0x16, 0x23, 0x0F, 0x23, 0x27, 0x03, 0x12, 0x20, 0x2F, 0x0D, 0x45,
	0x11, 0x2E, 0x3B, 0x0C, 0x3F, 0x52, 0x2E, 0x05, 0x15, 0x0A, 0x3A, 0x76,
	0x55, 0x51, 0x2F, 0x1F, 0x01, 0x3B, 0x11, 0x34, 0x38, 0x72, 0x59, 0x18,
	0x07, 0x39, 0x38, 0x02, 0x17, 0x2C, 0x2A, 0x08, 0x0F, 0x54, 0x17, 0x0E,
	0x09, 0x1B, 0x20, 0x38, 0x0F, 0x30, 0x14, 0x00, 0x2D, 0x5B, 0x18, 0x34,
	0x18, 0x24, 0x39, 0x7A, 0x05, 0x12, 0x0D, 0x40, 0x12, 0x22, 0x23, 0x26,
	0x0C, 0x13, 0x20, 0x2B, 0x1A, 0x1D, 0x34, 0x55, 0x37, 0x1E, 0x0F, 0x24,
	0x26, 0x52, 0x01, 0x25, 0x69, 0x3D, 0x36, 0x17, 0x53, 0x13, 0x02, 0x10,
	0x5C, 0x07, 0x03, 0x1C, 0x18, 0x02, 0x44, 0x1A, 0x19, 0x52, 0x3D, 0x08,
	0x2F, 0x20, 0x27, 0x3A, 0x5A, 0x0D, 0x3B, 0x12, 0x0F, 0x26, 0x0C, 0x3A,
	0x36, 0x28, 0x2A, 0x0C, 0x2F, 0x30, 0x36, 0x12, 0x38, 0x29, 0x3B, 0x23,
	0x5A, 0x73, 0x0B, 0x29, 0x5E, 0x22, 0x0C, 0x07, 0x10, 0x3D, 0x18, 0x70,
	0x5E, 0x0B, 0x25, 0x59, 0x11, 0x38, 0x13, 0x3A, 0x38, 0x73, 0x3D, 0x14,
	0x3C, 0x09, 0x13, 0x0F, 0x27, 0x39, 0x32, 0x0C, 0x2E, 0x2E, 0x28, 0x38,
	0x0F, 0x2F, 0x20, 0x41, 0x2C, 0x20, 0x1E, 0x10, 0x16, 0x5D, 0x20, 0x16,
	0x13, 0x3C, 0x5E, 0x74, 0x18, 0x2A, 0x19, 0x3F, 0x34, 0x3C, 0x02, 0x2F,
	0x33, 0x3B, 0x02, 0x16, 0x04, 0x1F, 0x03, 0x3A, 0x36, 0x1F, 0x1A, 0x2F,
	0x20, 0x19, 0x36, 0x1D, 0x30, 0x59, 0x36, 0x3B, 0x5A, 0x04, 0x19, 0x09,
	0x34, 0x1D, 0x1B, 0x04, 0x38, 0x23, 0x32, 0x71, 0x05, 0x05, 0x58, 0x03,
	0x15, 0x58, 0x39, 0x14, 0x28, 0x77, 0x2E, 0x24, 0x36, 0x5A, 0x0D, 0x14,
	0x2B, 0x5B, 0x1B, 0x37, 0x06, 0x35, 0x2A, 0x19, 0x24, 0x09, 0x2D, 0x22,
	0x5C, 0x38, 0x36, 0x23, 0x29, 0x18, 0x70, 0x54, 0x35, 0x1E, 0x0C, 0x73,
	0x28, 0x54, 0x27, 0x00, 0x11, 0x5E, 0x50, 0x16, 0x25, 0x7A, 0x2E, 0x02,
	0x39, 0x5B, 0x23, 0x18, 0x39, 0x38, 0x08, 0x0A, 0x0B, 0x22, 0x05, 0x59,
	0x2B, 0x1A, 0x28, 0x5C, 0x3E, 0x20, 0x58, 0x15, 0x3B, 0x08, 0x3A, 0x35,
	0x3B, 0x57, 0x3B, 0x14, 0x27, 0x00, 0x45, 0x5A, 0x13, 0x25, 0x51, 0x2C,
	0x32, 0x77, 0x26, 0x4E, 0x3C, 0x2C, 0x2F, 0x02, 0x11, 0x26, 0x04, 0x00,
	0x3C, 0x2F, 0x2F, 0x5B, 0x0C, 0x05, 0x2F, 0x0B, 0x3A, 0x28, 0x5F, 0x38,
	0x23, 0x1E, 0x33, 0x54, 0x2F, 0x5A, 0x0F, 0x25, 0x24, 0x2F, 0x3D, 0x52,
	0x7A, 0x19, 0x11, 0x39, 0x05, 0x09, 0x0F, 0x0E, 0x3B, 0x5E, 0x74, 0x3F,
	0x04, 0x04, 0x0E, 0x17, 0x06, 0x59, 0x45, 0x1E, 0x18, 0x55, 0x0D, 0x20,
	0x07, 0x0A, 0x5C, 0x2F, 0x34, 0x29, 0x26, 0x58, 0x33, 0x5A, 0x08, 0x03,
	0x08, 0x2B, 0x0D, 0x01, 0x76, 0x2A, 0x24, 0x01, 0x1E, 0x2B, 0x1C, 0x32,
	0x37, 0x2C, 0x30, 0x2F, 0x52, 0x25, 0x1F, 0x25, 0x02, 0x17, 0x00, 0x1E,
	0x13, 0x58, 0x2B, 0x59, 0x3E, 0x73, 0x1F, 0x0E, 0x24, 0x26, 0x2F, 0x1C,
	0x33, 0x0F, 0x28, 0x08, 0x3E, 0x06, 0x2B, 0x33, 0x3A, 0x01, 0x22, 0x0C,
	0x0D, 0x04, 0x3F, 0x34, 0x24, 0x12, 0x1A, 0x0D, 0x2C, 0x1A, 0x31, 0x09,
	0x23, 0x14, 0x23, 0x25, 0x17, 0x2F, 0x32, 0x19, 0x29, 0x2D, 0x1C, 0x29,
	0x23, 0x0F, 0x35, 0x5A, 0x1B, 0x04, 0x04, 0x70, 0x0B, 0x0B, 0x20, 0x20,
	0x77, 0x05, 0x58, 0x58, 0x5E, 0x0B, 0x5E, 0x03, 0x0C, 0x0D, 0x0E, 0x3C,
	0x0E, 0x09, 0x0E, 0x23, 0x5F, 0x0A, 0x05, 0x08, 0x27, 0x5D, 0x16, 0x01,
	0x0E, 0x3B, 0x5C, 0x16, 0x59, 0x29, 0x36, 0x5D, 0x16, 0x2F, 0x3A, 0x0A,
	0x0D, 0x39, 0x3F, 0x28, 0x33, 0x55, 0x09, 0x0A, 0x19, 0x04, 0x2A, 0x15,
	0x1D, 0x18, 0x6D, 0x01, 0x03, 0x14, 0x3F, 0x1B, 0x04, 0x17, 0x5C, 0x3A,
	0x14, 0x38, 0x58, 0x3D, 0x11, 0x35, 0x01, 0x14, 0x09, 0x5E, 0x25, 0x24,
	0x00, 0x1F, 0x40, 0x2E, 0x1C, 0x0C, 0x09, 0x23, 0x31, 0x0F, 0x23, 0x29,
	0x0C, 0x3A, 0x06, 0x2B, 0x1C, 0x20, 0x27, 0x27, 0x0C, 0x08, 0x3E, 0x04,
	0x3C, 0x28, 0x05, 0x0E, 0x71, 0x3E, 0x0E, 0x3F, 0x0F, 0x13, 0x28, 0x08,
	0x16, 0x1E, 0x09, 0x16, 0x20, 0x34, 0x25, 0x70, 0x5F, 0x06, 0x3F, 0x0A,
	0x33, 0x08, 0x04, 0x2F, 0x38, 0x0E, 0x3F, 0x4A, 0x2C, 0x31, 0x1A, 0x2E,
	0x30, 0x1D, 0x5E, 0x2F, 0x3B, 0x32, 0x5C, 0x5F, 0x04, 0x5D, 0x26, 0x22,
	0x1D, 0x72, 0x1C, 0x2A, 0x34, 0x02, 0x76, 0x23, 0x1B, 0x00, 0x44, 0x05,
	0x25, 0x27, 0x05, 0x24, 0x04, 0x36, 0x58, 0x18, 0x07, 0x73, 0x34, 0x33,
	0x45, 0x40, 0x32, 0x59, 0x50, 0x3D, 0x25, 0x10, 0x54, 0x12, 0x19, 0x52,
	0x30, 0x14, 0x26, 0x0B, 0x1F, 0x25, 0x1B, 0x37, 0x2C, 0x5D, 0x0C, 0x3B,
	0x25, 0x37, 0x27, 0x24, 0x26, 0x36, 0x0A, 0x3A, 0x3A, 0x5F, 0x3B, 0x03,
	0x3A, 0x0F, 0x1A, 0x17, 0x37, 0x26, 0x37, 0x34, 0x34, 0x56, 0x1F, 0x12,
	0x3D, 0x02, 0x18, 0x3A, 0x72, 0x01, 0x26, 0x0D, 0x38, 0x29, 0x43, 0x24,
	0x57, 0x5B, 0x0E, 0x29, 0x08, 0x5B, 0x11, 0x08, 0x24, 0x2D, 0x3C, 0x08,
	0x31, 0x05, 0x38, 0x18, 0x2F, 0x13, 0x28, 0x0C, 0x39, 0x1A, 0x0F, 0x38,
	0x4E, 0x08, 0x18, 0x0F, 0x07, 0x11, 0x16, 0x31, 0x00, 0x0D, 0x37, 0x2B,
	0x58, 0x15, 0x2A, 0x33, 0x18, 0x00, 0x23, 0x3F, 0x2B, 0x17, 0x0A, 0x05,
	0x35, 0x36, 0x1B, 0x52, 0x3B, 0x14, 0x0E, 0x2A, 0x33, 0x7B, 0x29, 0x13,
	0x58, 0x0C, 0x0B, 0x55, 0x30, 0x17, 0x03, 0x03, 0x28, 0x06, 0x38, 0x0D,
	0x07, 0x23, 0x39, 0x1E, 0x33, 0x0A, 0x2E, 0x2D, 0x3E, 0x2F, 0x6D, 0x06,
	0x4A, 0x5D, 0x22, 0x29, 0x0E, 0x51, 0x04, 0x32, 0x6D, 0x27, 0x36, 0x3B,
	0x38, 0x13, 0x21, 0x11, 0x1D, 0x1C, 0x25, 0x27, 0x23, 0x1D, 0x40, 0x27,
	0x1D, 0x2E, 0x28, 0x05, 0x08, 0x5F, 0x28, 0x29, 0x29, 0x07, 0x1C, 0x32,
	0x17, 0x38, 0x74, 0x39, 0x2C, 0x2D, 0x29, 0x0A, 0x1D, 0x10, 0x19, 0x11,
	0x32, 0x5A, 0x03, 0x01, 0x23, 0x1A, 0x07, 0x53, 0x24, 0x0F, 0x7B, 0x1F,
	0x2B, 0x3C, 0x1F, 0x70, 0x1C, 0x33, 0x05, 0x23, 0x2E, 0x25, 0x04, 0x5E,
	0x24, 0x24, 0x01, 0x08, 0x07, 0x08, 0x0B, 0x3E, 0x0F, 0x56, 0x59, 0x20,
	0x02, 0x53, 0x45, 0x19, 0x38, 0x2E, 0x58, 0x3E, 0x28, 0x3B, 0x5F, 0x51,
	0x17, 0x18, 0x6D, 0x24, 0x31, 0x5C, 0x24, 0x29, 0x0E, 0x0A, 0x00, 0x21,
	0x29, 0x29, 0x13, 0x45, 0x00, 0x2C, 0x27, 0x56, 0x23, 0x18, 0x18, 0x1F,
	0x34, 0x5E, 0x3F, 0x38, 0x0F, 0x0F, 0x3A, 0x04, 0x18, 0x22, 0x04, 0x25,
	0x21, 0x76, 0x58, 0x22, 0x20, 0x12, 0x30, 0x28, 0x27, 0x08, 0x38, 0x30,
	0x25, 0x2D, 0x19, 0x24, 0x26, 0x2D, 0x02, 0x1B, 0x5F, 0x7B, 0x47, 0x05,
	0x37, 0x20, 0x34, 0x0E, 0x27, 0x38, 0x12, 0x0F, 0x54, 0x2D, 0x01, 0x31,
	0x06, 0x21, 0x2F, 0x24, 0x5B, 0x08, 0x00, 0x50, 0x21, 0x0A, 0x6D, 0x28,
	0x53, 0x3C, 0x1D, 0x0A, 0x5F, 0x0E, 0x09, 0x27, 0x21, 0x2A, 0x07, 0x0F,
	0x2C, 0x09, 0x2F, 0x2D, 0x05, 0x2C, 0x2C, 0x2A, 0x22, 0x34, 0x5E, 0x38,
	0x1D, 0x03, 0x1F, 0x53, 0x00, 0x21, 0x06, 0x3B, 0x31, 0x30, 0x54, 0x28,
	0x3E, 0x09, 0x28, 0x15, 0x25, 0x09, 0x27, 0x73, 0x5A, 0x37, 0x0D, 0x28,
	0x73, 0x1F, 0x19, 0x0D, 0x3B, 0x32, 0x3C, 0x36, 0x1D, 0x00, 0x07, 0x03,
	0x2D, 0x22, 0x26, 0x37, 0x14, 0x19, 0x2B, 0x33, 0x03, 0x01, 0x2B, 0x38,
	0x2D, 0x33, 0x3F, 0x09, 0x3C, 0x08, 0x28, 0x2E, 0x51, 0x5A, 0x13, 0x27,
	0x3C, 0x25, 0x3F, 0x19, 0x7A, 0x58, 0x26, 0x04, 0x1B, 0x0B, 0x08, 0x2C,
	0x3D, 0x01, 0x0C, 0x28, 0x27, 0x28, 0x0F, 0x0E, 0x15, 0x29, 0x03, 0x59,
	0x01, 0x20, 0x18, 0x5C, 0x31, 0x06, 0x34, 0x53, 0x08, 0x3C, 0x26, 0x59,
	0x25, 0x3E, 0x5D, 0x11, 0x26, 0x32, 0x57, 0x5E, 0x01, 0x55, 0x28, 0x05,
	0x2C, 0x0E, 0x5F, 0x12, 0x06, 0x5A, 0x1B, 0x07, 0x35, 0x2F, 0x40, 0x18,
	0x1E, 0x0A, 0x2B, 0x00, 0x2B, 0x1D, 0x50, 0x2A, 0x08, 0x0F, 0x5D, 0x04,
	0x1F, 0x5F, 0x72, 0x0F, 0x33, 0x14, 0x18, 0x11, 0x3E, 0x58, 0x1A, 0x02,
	0x2F, 0x22, 0x29, 0x3A, 0x24, 0x69, 0x0D, 0x51, 0x0B, 0x3B, 0x69, 0x5A,
	0x0C, 0x0A, 0x24, 0x11, 0x14, 0x06, 0x19, 0x39, 0x01, 0x1F, 0x13, 0x2B,
	0x29, 0x16, 0x3E, 0x00, 0x0D, 0x08, 0x15, 0x3D, 0x23, 0x45, 0x53, 0x24,
	0x54, 0x15, 0x07, 0x3F, 0x06, 0x5C, 0x2D, 0x06, 0x1B, 0x03, 0x3E, 0x39,
	0x36, 0x03, 0x30, 0x23, 0x55, 0x16, 0x40, 0x2C, 0x03, 0x28, 0x45, 0x0D,
	0x13, 0x18, 0x36, 0x08, 0x09, 0x03, 0x1D, 0x19, 0x2F, 0x5F, 0x2F, 0x3A,
	0x2D, 0x19, 0x03, 0x12, 0x24, 0x56, 0x27, 0x24, 0x34, 0x1A, 0x34, 0x2A,
	0x23, 0x2B, 0x5E, 0x04, 0x00, 0x07, 0x03, 0x23, 0x24, 0x45, 0x5F, 0x31,
	0x36, 0x52, 0x04, 0x0C, 0x0C, 0x0E, 0x03, 0x0A, 0x2A, 0x0D, 0x06, 0x03,
	0x5B, 0x5B, 0x08, 0x22, 0x26, 0x34, 0x1A, 0x18, 0x01, 0x18, 0x39, 0x5F,
	0x09, 0x1B, 0x0B, 0x14, 0x01, 0x01, 0x0F, 0x09, 0x24, 0x59, 0x16, 0x15,
	0x28, 0x1E, 0x39, 0x03, 0x25, 0x52, 0x0B, 0x44, 0x13, 0x0D, 0x0C, 0x03,
	0x1B, 0x2A, 0x1A, 0x28, 0x41, 0x0C, 0x37, 0x36, 0x11, 0x06, 0x23, 0x76,
	0x47, 0x31, 0x18, 0x24, 0x31, 0x27, 0x13, 0x3A, 0x3A, 0x27, 0x26, 0x2F,
	0x41, 0x5F, 0x25, 0x24, 0x0A, 0x2D, 0x2C, 0x1B, 0x1B, 0x39, 0x5A, 0x5B,
	0x2F, 0x1B, 0x24, 0x0D, 0x22, 0x26, 0x3C, 0x05, 0x24, 0x58, 0x2A, 0x22,
	0x24, 0x16, 0x3F, 0x21, 0x34, 0x0C, 0x1F, 0x02, 0x0B, 0x2B, 0x51, 0x01,
	0x04, 0x0D, 0x23, 0x2F, 0x3B, 0x2D, 0x20, 0x15, 0x32, 0x03, 0x05, 0x77,
	0x23, 0x2D, 0x41, 0x08, 0x18, 0x26, 0x0E, 0x5D, 0x11, 0x03, 0x01, 0x1B,
	0x0D, 0x1C, 0x04, 0x54, 0x09, 0x26, 0x27, 0x29, 0x1A, 0x30, 0x07, 0x31,
	0x70, 0x07, 0x57, 0x3A, 0x0A, 0x16, 0x3F, 0x08, 0x05, 0x06, 0x7A, 0x04,
	0x0F, 0x58, 0x2A, 0x18, 0x01, 0x54, 0x57, 0x21, 0x01, 0x2F, 0x34, 0x5D,
	0x03, 0x07, 0x1B, 0x2B, 0x5E, 0x2E, 0x0F, 0x00, 0x03, 0x5A, 0x22, 0x08,
	0x39, 0x11, 0x5D, 0x04, 0x00, 0x3C, 0x2E, 0x5B, 0x06, 0x14, 0x22, 0x50,
	0x00, 0x24, 0x06, 0x26, 0x20, 0x09, 0x22, 0x09, 0x43, 0x0A, 0x1C, 0x12,
	0x32, 0x59, 0x2B, 0x08, 0x19, 0x0E, 0x07, 0x37, 0x09, 0x52, 0x69, 0x06,
	0x39, 0x02, 0x0D, 0x08, 0x1A, 0x19, 0x20, 0x40, 0x6D, 0x1B, 0x29, 0x0B,
	0x09, 0x70, 0x2B, 0x53, 0x09, 0x19, 0x35, 0x09, 0x05, 0x23, 0x2E, 0x04,
	0x2F, 0x52, 0x26, 0x0C, 0x15, 0x5D, 0x20, 0x0A, 0x11, 0x00, 0x3A, 0x05,
	0x24, 0x5B, 0x0D, 0x23, 0x34, 0x3A, 0x03, 0x11, 0x26, 0x20, 0x27, 0x0A,
	0x7B, 0x55, 0x37, 0x39, 0x1E, 0x1B, 0x01, 0x36, 0x45, 0x32, 0x36, 0x01,
	0x06, 0x1B, 0x13, 0x25, 0x07, 0x24, 0x0A, 0x33, 0x29, 0x5B, 0x54, 0x57,
	0x3F, 0x77, 0x3E, 0x4A, 0x5F, 0x3E, 0x34, 0x23, 0x0A, 0x2C, 0x04, 0x33,
	0x39, 0x37, 0x18, 0x40, 0x76, 0x28, 0x2A, 0x20, 0x1D, 0x77, 0x2B, 0x18,
	0x26, 0x0A, 0x35, 0x1C, 0x19, 0x0B, 0x5C, 0x0F, 0x00, 0x07, 0x16, 0x52,
	0x75, 0x5E, 0x15, 0x04, 0x03, 0x76, 0x5A, 0x09, 0x1B, 0x5B, 0x09, 0x0B,
	0x3B, 0x45, 0x1E, 0x09, 0x36, 0x2E, 0x1F, 0x22, 0x2C, 0x5F, 0x04, 0x57,
	0x05, 0x37, 0x28, 0x0E, 0x3E, 0x22, 0x2E, 0x22, 0x2F, 0x25, 0x0C, 0x73,
	0x2D, 0x54, 0x04, 0x07, 0x28, 0x5F, 0x55, 0x03, 0x0D, 0x0E, 0x08, 0x23,
	0x3D, 0x13, 0x75, 0x0A, 0x50, 0x28, 0x5F, 0x30, 0x08, 0x36, 0x14, 0x3D,
	0x08, 0x07, 0x27, 0x5B, 0x0F, 0x11, 0x0B, 0x11, 0x19, 0x08, 0x23, 0x26,
	0x4A, 0x2A, 0x1F, 0x71, 0x2D, 0x27, 0x1B, 0x0C, 0x2A, 0x2B, 0x20, 0x0C,
	0x59, 0x25, 0x3C, 0x0C, 0x39, 0x3B, 0x3B, 0x47, 0x27, 0x3C, 0x2D, 0x29,
	0x29, 0x30, 0x00, 0x1E, 0x07, 0x0F, 0x0C, 0x09, 0x03, 0x1B, 0x05, 0x06,
	0x04, 0x26, 0x03, 0x0B, 0x22, 0x04, 0x59, 0x69, 0x59, 0x4E, 0x01, 0x2A,
	0x17, 0x07, 0x0D, 0x17, 0x25, 0x7B, 0x3E, 0x04, 0x2F, 0x20, 0x10, 0x35,
	0x54, 0x1D, 0x5E, 0x75, 0x15, 0x56, 0x20, 0x52, 0x2D, 0x02, 0x05, 0x0F,
	0x3C, 0x34, 0x03, 0x2A, 0x57, 0x24, 0x2D, 0x0F, 0x27, 0x14, 0x40, 0x1A,
	0x1A, 0x2A, 0x0F, 0x27, 0x75, 0x38, 0x08, 0x0D, 0x18, 0x20, 0x2F, 0x2C,
	0x01, 0x27, 0x31, 0x38, 0x18, 0x07, 0x0A, 0x71, 0x58, 0x35, 0x04, 0x2C,
	0x32, 0x1C, 0x0A, 0x02, 0x38, 0x06, 0x0E, 0x0B, 0x2B, 0x0C, 0x76, 0x2B,
	0x2F, 0x00, 0x33, 0x13, 0x16, 0x11, 0x16, 0x39, 0x1B, 0x2E, 0x39, 0x17,
	0x33, 0x7B, 0x5A, 0x0B, 0x5B, 0x12, 0x10, 0x36, 0x16, 0x00, 0x3E, 0x37,
	0x3F, 0x23, 0x1D, 0x2F, 0x13, 0x20, 0x53, 0x1A, 0x20, 0x7B, 0x3D, 0x09,
	0x21, 0x32, 0x7B, 0x5D, 0x2B, 0x05, 0x23, 0x09, 0x22, 0x31, 0x27, 0x5A,
	0x6D, 0x0E, 0x09, 0x2B, 0x1B, 0x3A, 0x2B, 0x3B, 0x5F, 0x01, 0x6D, 0x2D,
	0x00, 0x41, 0x3D, 0x0F, 0x59, 0x25, 0x5D, 0x20, 0x01, 0x2A, 0x25, 0x58,
	0x3F, 0x0B, 0x43, 0x07, 0x01, 0x12, 0x27, 0x35, 0x04, 0x37, 0x59, 0x34,
	0x0D, 0x02, 0x3E, 0x22, 0x3A, 0x36, 0x57, 0x14, 0x39, 0x05, 0x0B, 0x59,
	0x3D, 0x5F, 0x10, 0x2A, 0x2C, 0x09, 0x1E, 0x7B, 0x2F, 0x15, 0x27, 0x20,
	0x33, 0x2A, 0x12, 0x18, 0x44, 0x77, 0x1B, 0x24, 0x3B, 0x0C, 0x0E, 0x09,
	0x29, 0x56, 0x2A, 0x6D, 0x35, 0x57, 0x29, 0x3F, 0x24, 0x23, 0x16, 0x39,
	0x13, 0x71, 0x2D, 0x03, 0x18, 0x2F, 0x3B, 0x2D, 0x31, 0x39, 0x27, 0x0D,
	0x26, 0x29, 0x3B, 0x12, 0x15, 0x23, 0x17, 0x26, 0x03, 0x11, 0x0F, 0x0D,
	0x26, 0x23, 0x70, 0x55, 0x51, 0x25, 0x18, 0x0A, 0x20, 0x2F, 0x24, 0x26,
	0x2A, 0x07, 0x4E, 0x3F, 0x12, 0x33, 0x09, 0x15, 0x45, 0x07, 0x28, 0x55,
	0x29, 0x00, 0x0C, 0x2F, 0x1F, 0x27, 0x5F, 0x21, 0x1A, 0x1D, 0x15, 0x16,
	0x33, 0x2F, 0x2F, 0x06, 0x19, 0x2E, 0x07, 0x5B, 0x55, 0x59, 0x44, 0x32,
	0x35, 0x2F, 0x26, 0x44, 0x0E, 0x0A, 0x59, 0x28, 0x08, 0x7A, 0x43, 0x2A,
	0x45, 0x28, 0x69, 0x03, 0x59, 0x04, 0x0A, 0x6D, 0x5E, 0x0C, 0x39, 0x3E,
	0x74, 0x47, 0x0E, 0x1F, 0x09, 0x32, 0x3E, 0x0C, 0x5B, 0x2F, 0x2E, 0x2D,
	0x11, 0x0B, 0x3F, 0x75, 0x3D, 0x4A, 0x0B, 0x01, 0x04, 0x25, 0x2F, 0x3E,
	0x39, 0x01, 0x34, 0x07, 0x2C, 0x2A, 0x2F, 0x02, 0x35, 0x05, 0x22, 0x2C,
	0x19, 0x0C, 0x1F, 0x59, 0x69, 0x24, 0x36, 0x59, 0x13, 0x15, 0x5B, 0x19,
	0x45, 0x1E, 0x76, 0x18, 0x2F, 0x16, 0x08, 0x2D, 0x43, 0x2E, 0x0F, 0x3F,
	0x16, 0x2D, 0x58, 0x02, 0x5C, 0x06, 0x5E, 0x24, 0x0B, 0x1B, 0x2C, 0x3C,
	0x0C, 0x3D, 0x18, 0x32, 0x14, 0x08, 0x5E, 0x05, 0x3B, 0x38, 0x58, 0x06,
	0x03, 0x26, 0x00, 0x20, 0x0C, 0x5A, 0x20, 0x34, 0x56, 0x1B, 0x2E, 0x71,
	0x27, 0x24, 0x02, 0x40, 0x0F, 0x2F, 0x25, 0x39, 0x28, 0x30, 0x21, 0x4A,
	0x3F, 0x24, 0x3A, 0x38, 0x0B, 0x2C, 0x52, 0x01, 0x07, 0x33, 0x1D, 0x3E,
	0x25, 0x55, 0x59, 0x1B, 0x0D, 0x04, 0x0B, 0x15, 0x14, 0x3B, 0x08, 0x3F,
	0x38, 0x1B, 0x1B, 0x30, 0x5E, 0x2A, 0x2D, 0x38, 0x69, 0x04, 0x16, 0x45,
	0x1C, 0x01, 0x03, 0x11, 0x14, 0x3B, 0x1B, 0x2A, 0x2D, 0x5C, 0x3B, 0x38,
	0x19, 0x0D, 0x5B, 0x21, 0x15, 0x01, 0x4E, 0x5D, 0x19, 0x0A, 0x34, 0x04,
	0x0F, 0x58, 0x12, 0x59, 0x59, 0x00, 0x2E, 0x15, 0x2B, 0x37, 0x3B, 0x59,
	0x11, 0x5F, 0x39, 0x16, 0x3D, 0x03, 0x02, 0x54, 0x41, 0x20, 0x76, 0x07,
	0x34, 0x0B, 0x0E, 0x12, 0x06, 0x06, 0x27, 0x0C, 0x01, 0x22, 0x25, 0x1C,
	0x08, 0x2D, 0x3C, 0x32, 0x2C, 0x5D, 0x30, 0x39, 0x2E, 0x02, 0x09, 0x0E,
	0x01, 0x50, 0x14, 0x5C, 0x2A, 0x5C, 0x31, 0x00, 0x5D, 0x76, 0x03, 0x12,
	0x5C, 0x22, 0x35, 0x22, 0x33, 0x2C, 0x40, 0x7A, 0x24, 0x38, 0x3B, 0x29,
	0x04, 0x02, 0x4E, 0x3E, 0x20, 0x2E, 0x0F, 0x19, 0x5E, 0x04, 0x08, 0x47,
	0x10, 0x29, 0x13, 0x35, 0x3E, 0x57, 0x00, 0x22, 0x2D, 0x5E, 0x22, 0x2C,
	0x31, 0x0B, 0x5E, 0x14, 0x1D, 0x2D, 0x09, 0x1B, 0x2F, 0x09, 0x1A, 0x03,
	0x0E, 0x23, 0x57, 0x3C, 0x2B, 0x0E, 0x55, 0x14, 0x3F, 0x21, 0x3F, 0x37,
	0x20, 0x58, 0x37, 0x1B, 0x0F, 0x1A, 0x3B, 0x73, 0x55, 0x36, 0x36, 0x33,
	0x37, 0x04, 0x11, 0x36, 0x02, 0x74, 0x5A, 0x59, 0x1A, 0x58, 0x0A, 0x1E,
	0x30, 0x00, 0x02, 0x73, 0x1E, 0x2C, 0x2F, 0x19, 0x77, 0x1F, 0x2F, 0x1F,
	0x59, 0x29, 0x59, 0x34, 0x07, 0x5D, 0x03, 0x3A, 0x36, 0x41, 0x1C, 0x03,
	0x1A, 0x23, 0x08, 0x3A, 0x0B, 0x1D, 0x1B, 0x5E, 0x00, 0x71, 0x29, 0x12,
	0x04, 0x20, 0x35, 0x2E, 0x23, 0x02, 0x52, 0x11, 0x14, 0x36, 0x39, 0x03,
	0x00, 0x24, 0x20, 0x08, 0x22, 0x7A, 0x0E, 0x53, 0x0F, 0x3E, 0x2B, 0x2D,
	0x19, 0x34, 0x00, 0x0B, 0x23, 0x2B, 0x09, 0x5E, 0x05, 0x1D, 0x0B, 0x1A,
	0x32, 0x34, 0x3F, 0x20, 0x25, 0x3F, 0x29, 0x3C, 0x2F, 0x18, 0x2D, 0x2D,
	0x1D, 0x18, 0x1C, 0x53, 0x0B, 0x1B, 0x08, 0x05, 0x3B, 0x04, 0x16, 0x34,
	0x25, 0x39, 0x27, 0x20, 0x52, 0x04, 0x2E, 0x74, 0x39, 0x35, 0x0C, 0x0F,
	0x27, 0x1C, 0x28, 0x56, 0x38, 0x37, 0x23, 0x19, 0x34, 0x0D, 0x2C, 0x18,
	0x12, 0x1B, 0x19, 0x75, 0x2B, 0x3B, 0x25, 0x3F, 0x03, 0x1D, 0x25, 0x20,
	0x2F, 0x73, 0x03, 0x56, 0x23, 0x3A, 0x32, 0x0D, 0x53, 0x5D, 0x2E, 0x09,
	0x47, 0x12, 0x38, 0x06, 0x0E, 0x03, 0x30, 0x58, 0x1C, 0x18, 0x55, 0x2A,
	0x16, 0x31, 0x0B, 0x54, 0x24, 0x41, 0x11, 0x01, 0x59, 0x08, 0x0C, 0x58,
	0x2A, 0x07, 0x2A, 0x5F, 0x3C, 0x05, 0x0B, 0x3B, 0x28, 0x01, 0x0E, 0x55,
	0x04, 0x3F, 0x3F, 0x77, 0x55, 0x29, 0x0C, 0x23, 0x07, 0x05, 0x0B, 0x57,
	0x21, 0x38, 0x3D, 0x05, 0x08, 0x28, 0x2C, 0x21, 0x1B, 0x5D, 0x22, 0x2A,
	0x59, 0x05, 0x2B, 0x3C, 0x7A, 0x07, 0x12, 0x5B, 0x53, 0x08, 0x2A, 0x33,
	0x2C, 0x1E, 0x38, 0x1F, 0x08, 0x2A, 0x2F, 0x75, 0x23, 0x09, 0x25, 0x13,
	0x36, 0x58, 0x2E, 0x1A, 0x1E, 0x74, 0x08, 0x2B, 0x1A, 0x2C, 0x35, 0x38,
	0x39, 0x21, 0x0F, 0x28, 0x3D, 0x12, 0x05, 0x1B, 0x71, 0x23, 0x08, 0x0D,
	0x53, 0x32, 0x1B, 0x13, 0x59, 0x11, 0x69, 0x34, 0x20, 0x24, 0x2A, 0x03,
	0x2E, 0x2D, 0x20, 0x3B, 0x74, 0x2A, 0x29, 0x03, 0x5D, 0x0E, 0x05, 0x4A,
	0x3E, 0x0C, 0x23, 0x19, 0x19, 0x17, 0x2E, 0x00, 0x22, 0x2C, 0x38, 0x0A,
	0x06, 0x19, 0x26, 0x02, 0x1C, 0x13, 0x22, 0x3B, 0x38, 0x25, 0x04, 0x3E,
	0x0F, 0x07, 0x25, 0x35, 0x23, 0x2E, 0x45, 0x28, 0x25, 0x38, 0x56, 0x39,
	0x04, 0x25, 0x5E, 0x51, 0x3E, 0x1C, 0x35, 0x5C, 0x38, 0x16, 0x3A, 0x28,
	0x43, 0x52, 0x3D, 0x5A, 0x05, 0x58, 0x52, 0x5C, 0x24, 0x2A, 0x15, 0x15,
	0x09, 0x1D, 0x35, 0x09, 0x54, 0x27, 0x20, 0x2C, 0x01, 0x0F, 0x04, 0x0D,
	0x0C, 0x05, 0x09, 0x5D, 0x27, 0x29, 0x5B, 0x0E, 0x59, 0x21, 0x76, 0x07,
	0x23, 0x20, 0x33, 0x30, 0x3D, 0x3B, 0x0D, 0x00, 0x04, 0x58, 0x36, 0x01,
	0x38, 0x71, 0x5F, 0x0A, 0x2C, 0x24, 0x2F, 0x0A, 0x14, 0x3F, 0x2A, 0x2B,
	0x27, 0x27, 0x34, 0x06, 0x01, 0x16, 0x04, 0x5D, 0x18, 0x32, 0x34, 0x06,
	0x08, 0x0E, 0x0B, 0x1B, 0x06, 0x59, 0x0E, 0x32, 0x2A, 0x02, 0x1A, 0x39,
	0x35, 0x15, 0x36, 0x1A, 0x5A, 0x0A, 0x1F, 0x4E, 0x25, 0x3B, 0x76, 0x59,
	0x27, 0x28, 0x0F, 0x0E, 0x3B, 0x19, 0x05, 0x18, 0x16, 0x3A, 0x14, 0x04,
	0x39, 0x1A, 0x06, 0x09, 0x2C, 0x23, 0x08, 0x43, 0x36, 0x2F, 0x2F, 0x34,
	0x27, 0x27, 0x09, 0x0A, 0x76, 0x1B, 0x59, 0x00, 0x12, 0x0C, 0x23, 0x16,
	0x1E, 0x03, 0x2F, 0x0E, 0x05, 0x57, 0x0D, 0x13, 0x5C, 0x0F, 0x06, 0x27,
	0x33, 0x35, 0x23, 0x1D, 0x1E, 0x2A, 0x25, 0x1B, 0x0A, 0x38, 0x00, 0x1F,
	0x34, 0x5F, 0x24, 0x28, 0x0B, 0x58, 0x26, 0x3C, 0x33, 0x5B, 0x2A, 0x56,
	0x02, 0x26, 0x1B, 0x0F, 0x1C, 0x3E, 0x27, 0x29, 0x54, 0x58, 0x58, 0x0B,
	0x5E, 0x56, 0x29, 0x01, 0x08, 0x5A, 0x23, 0x37, 0x53, 0x0F, 0x5D, 0x38,
	0x0B, 0x04, 0x38, 0x0D, 0x35, 0x5D, 0x05, 0x71, 0x22, 0x05, 0x21, 0x20,
	0x7B, 0x21, 0x00, 0x03, 0x44, 0x03, 0x24, 0x30, 0x3E, 0x11, 0x1B, 0x2E,
	0x2B, 0x17, 0x1D, 0x18, 0x06, 0x1B, 0x16, 0x2E, 0x0E, 0x27, 0x0D, 0x5A,
	0x39, 0x29, 0x25, 0x0C, 0x23, 0x0D, 0x2B, 0x29, 0x00, 0x3E, 0x05, 0x04,
	0x0F, 0x3B, 0x05, 0x04, 0x33, 0x54, 0x27, 0x0B, 0x08, 0x1A, 0x16, 0x25,
	0x3B, 0x1E, 0x71, 0x03, 0x2D, 0x5F, 0x04, 0x15, 0x25, 0x31, 0x20, 0x1C,
	0x00, 0x03, 0x0F, 0x1C, 0x39, 0x2C, 0x3E, 0x1B, 0x25, 0x1A, 0x27, 0x5A,
	0x0D, 0x1B, 0x19, 0x0B, 0x3F, 0x16, 0x18, 0x3A, 0x2F, 0x5E, 0x27, 0x0A,
	0x2F, 0x33, 0x25, 0x38, 0x06, 0x20, 0x14, 0x5A, 0x1B, 0x59, 0x07, 0x74,
	0x3A, 0x22, 0x06, 0x2A, 0x33, 0x29, 0x06, 0x5E, 0x3A, 0x23, 0x1D, 0x31,
	0x1E, 0x0E, 0x10, 0x2A, 0x50, 0x25, 0x19, 0x01, 0x28, 0x53, 0x5E, 0x06,
	0x15, 0x09, 0x24, 0x5E, 0x29, 0x69, 0x43, 0x32, 0x45, 0x02, 0x31, 0x2A,
	0x00, 0x3F, 0x1F, 0x2B, 0x0D, 0x22, 0x37, 0x40, 0x20, 0x22, 0x09, 0x09,
	0x19, 0x27, 0x21, 0x10, 0x3B, 0x0A, 0x75, 0x3B, 0x2E, 0x07, 0x44, 0x23,
	0x27, 0x02, 0x02, 0x12, 0x0B, 0x1E, 0x34, 0x17, 0x03, 0x38, 0x5D, 0x2A,
	0x39, 0x2E, 0x05, 0x3D, 0x28, 0x05, 0x00, 0x2C, 0x2D, 0x17, 0x56, 0x29,
	0x11, 0x2B, 0x35, 0x59, 0x2A, 0x37, 0x23, 0x3B, 0x07, 0x5D, 0x23, 0x2D,
	0x59, 0x02, 0x00, 0x3A, 0x35, 0x4A, 0x5C, 0x0D, 0x0B, 0x22, 0x3B, 0x56,
	0x1C, 0x17, 0x5F, 0x19, 0x57, 0x19, 0x33, 0x07, 0x52, 0x2F, 0x02, 0x2F,
	0x35, 0x37, 0x45, 0x0C, 0x27, 0x3B, 0x20, 0x24, 0x0C, 0x34, 0x18, 0x39,
	0x5B, 0x2F, 0x26, 0x15, 0x25, 0x36, 0x2F, 0x26, 0x15, 0x4E, 0x57, 0x00,
	0x1B, 0x20, 0x28, 0x06, 0x04, 0x7B, 0x5E, 0x0D, 0x1F, 0x09, 0x2A, 0x3A,
	0x0B, 0x23, 0x33, 0x0D, 0x25, 0x33, 0x5A, 0x5D, 0x03, 0x20, 0x0B, 0x38,
	0x2C, 0x2B, 0x0B, 0x37, 0x3E, 0x2A, 0x34, 0x00, 0x04, 0x06, 0x03, 0x0D,
	0x0F, 0x59, 0x22, 0x53, 0x73, 0x3D, 0x4E, 0x56, 0x2D, 0x1A, 0x0B, 0x37,
	0x03, 0x2E, 0x08, 0x3B, 0x54, 0x05, 0x3E, 0x00, 0x22, 0x06, 0x1E, 0x18,
	0x0D, 0x1B, 0x37, 0x39, 0x0E, 0x73, 0x07, 0x35, 0x1C, 0x04, 0x11, 0x04,
	0x19, 0x00, 0x31, 0x08, 0x3C, 0x0B, 0x2C, 0x53, 0x13, 0x58, 0x50, 0x0A,
	0x38, 0x13, 0x3D, 0x04, 0x5B, 0x19, 0x2A, 0x34, 0x20, 0x1F, 0x58, 0x23,
	0x15, 0x57, 0x41, 0x5F, 0x25, 0x5B, 0x06, 0x0D, 0x27, 0x04, 0x2D, 0x2F,
	0x58, 0x5A, 0x25, 0x21, 0x05, 0x5C, 0x13, 0x2A, 0x16, 0x2F, 0x1B, 0x26,
	0x24, 0x05, 0x31, 0x1D, 0x1E, 0x06, 0x0A, 0x38, 0x41, 0x40, 0x04, 0x47,
	0x2F, 0x0C, 0x5F, 0x37, 0x1F, 0x0F, 0x5B, 0x29, 0x10, 0x05, 0x09, 0x04,
	0x2E, 0x28, 0x34, 0x0C, 0x2A, 0x03, 0x73, 0x34, 0x08, 0x08, 0x22, 0x1B,
	0x55, 0x20, 0x02, 0x1C, 0x18, 0x26, 0x0F, 0x16, 0x3D, 0x3A, 0x14, 0x25,
	0x0B, 0x0F, 0x2B, 0x43, 0x2E, 0x18, 0x2A, 0x29, 0x2D, 0x08, 0x1C, 0x24,
	0x2C, 0x5A, 0x22, 0x23, 0x26, 0x0C, 0x18, 0x06, 0x29, 0x2F, 0x0E, 0x14,
	0x35, 0x0B, 0x2A, 0x28, 0x2D, 0x0E, 0x07, 0x1C, 0x77, 0x5B, 0x58, 0x2B,
	0x2F, 0x27, 0x26, 0x10, 0x5E, 0x05, 0x14, 0x23, 0x55, 0x01, 0x5C, 0x0E,
	0x00, 0x26, 0x58, 0x1E, 0x25, 0x22, 0x0D, 0x41, 0x26, 0x31, 0x2A, 0x13,
	0x20, 0x08, 0x0C, 0x5C, 0x50, 0x25, 0x26, 0x35, 0x18, 0x06, 0x39, 0x0C,
	0x35, 0x1A, 0x12, 0x02, 0x1E, 0x1B, 0x54, 0x07, 0x2B, 0x19, 0x1B, 0x09,
	0x06, 0x0B, 0x0A, 0x14, 0x39, 0x36, 0x2A, 0x1B, 0x08, 0x5C, 0x26, 0x3D,
	0x33, 0x33, 0x1B, 0x02, 0x05, 0x32, 0x2B, 0x18, 0x53, 0x19, 0x2E, 0x71,
	0x5B, 0x0A, 0x36, 0x2C, 0x75, 0x23, 0x37, 0x41, 0x24, 0x24, 0x59, 0x31,
	0x5E, 0x27, 0x72, 0x3D, 0x0E, 0x3E, 0x18, 0x25, 0x3D, 0x22, 0x24, 0x04,
	0x2B, 0x1F, 0x07, 0x2A, 0x0E, 0x12, 0x05, 0x10, 0x3D, 0x38, 0x25, 0x2A,
	0x53, 0x3C, 0x13, 0x7B, 0x29, 0x12, 0x16, 0x13, 0x77, 0x1D, 0x08, 0x45,
	0x29, 0x32, 0x15, 0x0F, 0x36, 0x2E, 0x15, 0x58, 0x34, 0x2C, 0x1B, 0x3A,
	0x58, 0x08, 0x1C, 0x2C, 0x28, 0x2F, 0x2C, 0x27, 0x3A, 0x37, 0x23, 0x57,
	0x0C, 0x3F, 0x3A, 0x03, 0x00, 0x26, 0x25, 0x08, 0x3E, 0x4E, 0x5F, 0x12,
	0x05, 0x5E, 0x11, 0x3D, 0x11, 0x29, 0x09, 0x20, 0x22, 0x2D, 0x38, 0x24,
	0x18, 0x0D, 0x33, 0x37, 0x3C, 0x0A, 0x59, 0x02, 0x16, 0x0E, 0x18, 0x2B,
	0x0D, 0x35, 0x2A, 0x4E, 0x24, 0x0D, 0x03, 0x27, 0x31, 0x07, 0x5C, 0x2A,
	0x1C, 0x51, 0x28, 0x21, 0x27, 0x24, 0x12, 0x0D, 0x23, 0x77, 0x36, 0x10,
	0x3B, 0x09, 0x25, 0x2E, 0x25, 0x27, 0x04, 0x06, 0x2F, 0x3B, 0x2C, 0x12,
	0x08, 0x47, 0x3B, 0x04, 0x02, 0x2E, 0x3D, 0x0C, 0x2A, 0x1E, 0x0F, 0x02,
	0x30, 0x26, 0x5C, 0x3A, 0x3D, 0x26, 0x06, 0x05, 0x75, 0x05, 0x23, 0x23,
	0x5E, 0x25, 0x54, 0x23, 0x01, 0x22, 0x14, 0x34, 0x51, 0x20, 0x58, 0x04,
	0x34, 0x2C, 0x21, 0x07, 0x2E, 0x0A, 0x16, 0x38, 0x59, 0x73, 0x06, 0x38,
	0x3F, 0x31, 0x2B, 0x25, 0x0A, 0x1B, 0x40, 0x2F, 0x08, 0x3B, 0x2B, 0x0D,
	0x20, 0x58, 0x27, 0x3C, 0x05, 0x05, 0x07, 0x06, 0x3D, 0x5C, 0x07, 0x2A,
	0x36, 0x0F, 0x09, 0x01, 0x5F, 0x51, 0x1A, 0x2F, 0x0F, 0x25, 0x51, 0x06,
	0x32, 0x09, 0x00, 0x57, 0x58, 0x24, 0x71, 0x19, 0x16, 0x56, 0x0C, 0x37,
	0x28, 0x26, 0x3E, 0x3A, 0x31, 0x1F, 0x0A, 0x16, 0x3A, 0x3A, 0x47, 0x2A,
	0x0F, 0x3A, 0x13, 0x07, 0x20, 0x37, 0x5B, 0x29, 0x0B, 0x31, 0x3B, 0x20,
	0x2A, 0x21, 0x35, 0x05, 0x18, 0x2F, 0x16, 0x02, 0x07, 0x1C, 0x70, 0x04,
	0x56, 0x07, 0x44, 0x38, 0x22, 0x07, 0x2F, 0x11, 0x29, 0x2D, 0x1B, 0x2F,
	0x3A, 0x0A, 0x5C, 0x08, 0x0F, 0x03, 0x34, 0x16, 0x59, 0x00, 0x2E, 0x7B,
	0x5C, 0x56, 0x21, 0x21, 0x05, 0x0E, 0x13, 0x17, 0x1B, 0x2A, 0x59, 0x29,
	0x03, 0x0E, 0x13, 0x19, 0x28, 0x5C, 0x1D, 0x28, 0x5A, 0x16, 0x23, 0x53,
	0x7A, 0x1D, 0x36, 0x20, 0x40, 0x6D, 0x3F, 0x02, 0x36, 0x24, 0x1B, 0x43,
	0x0A, 0x24, 0x03, 0x26, 0x26, 0x08, 0x17, 0x1F, 0x04, 0x36, 0x39, 0x45,
	0x25, 0x21, 0x28, 0x19, 0x00, 0x3C, 0x21, 0x24, 0x58, 0x18, 0x3C, 0x06,
	0x09, 0x03, 0x28, 0x5A, 0x0D, 0x3E, 0x05, 0x3D, 0x29, 0x12, 0x0A, 0x31,
	0x05, 0x2F, 0x00, 0x1F, 0x3B, 0x25, 0x27, 0x38, 0x05, 0x2D, 0x2C, 0x5B,
	0x7B, 0x2A, 0x39, 0x1B, 0x1F, 0x1B, 0x26, 0x29, 0x09, 0x3C, 0x18, 0x0F,
	0x07, 0x02, 0x58, 0x70, 0x03, 0x04, 0x14, 0x3A, 0x2C, 0x22, 0x27, 0x36,
	0x29, 0x11, 0x54, 0x2F, 0x5C, 0x52, 0x2C, 0x27, 0x15, 0x37, 0x06, 0x37,
	0x3F, 0x14, 0x2C, 0x53, 0x24, 0x24, 0x07, 0x1D, 0x1D, 0x34, 0x20, 0x00,
	0x3C, 0x21, 0x18, 0x5A, 0x32, 0x5A, 0x1A, 0x2D, 0x55, 0x20, 0x14, 0x0F,
	0x29, 0x0B, 0x16, 0x1E, 0x20, 0x11, 0x15, 0x27, 0x2A, 0x13, 0x3A, 0x06,
	0x00, 0x1B, 0x3F, 0x18, 0x1B, 0x26, 0x5F, 0x44, 0x2A, 0x08, 0x59, 0x0B,
	0x00, 0x0B, 0x0F, 0x27, 0x03, 0x08, 0x27, 0x3C, 0x0A, 0x1E, 0x1D, 0x15,
	0x19, 0x05, 0x3F, 0x3F, 0x35, 0x04, 0x19, 0x45, 0x2F, 0x75, 0x59, 0x03,
	0x38, 0x2E, 0x26, 0x5F, 0x2C, 0x3B, 0x26, 0x14, 0x08, 0x07, 0x19, 0x24,
	0x27, 0x27, 0x51, 0x37, 0x0E, 0x14, 0x39, 0x12, 0x0A, 0x5D, 0x08, 0x47,
	0x09, 0x39, 0x3E, 0x28, 0x0F, 0x50, 0x5E, 0x40, 0x2C, 0x0E, 0x22, 0x1D,
	0x1E, 0x37, 0x58, 0x20, 0x3F, 0x20, 0x36, 0x24, 0x15, 0x03, 0x40, 0x2B,
	0x3C, 0x25, 0x27, 0x58, 0x21, 0x2D, 0x07, 0x07, 0x3B, 0x6D, 0x1B, 0x28,
	0x0C, 0x04, 0x75, 0x58, 0x20, 0x36, 0x01, 0x0E, 0x5C, 0x35, 0x06, 0x52,
	0x74, 0x55, 0x4E, 0x5A, 0x3E, 0x73, 0x08, 0x23, 0x02, 0x33, 0x6D, 0x00,
	0x35, 0x19, 0x3E, 0x69, 0x1B, 0x54, 0x09, 0x29, 0x2D, 0x2B, 0x56, 0x5D,
	0x02, 0x04, 0x18, 0x37, 0x20, 0x3D, 0x3B, 0x1A, 0x32, 0x29, 0x33, 0x77,
	0x1F, 0x09, 0x56, 0x3D, 0x05, 0x23, 0x27, 0x2A, 0x0D, 0x73, 0x2A, 0x17,
	0x06, 0x03, 0x3A, 0x5D, 0x0B, 0x0F, 0x24, 0x74, 0x2A, 0x3B, 0x3A, 0x07,
	0x2B, 0x5A, 0x55, 0x3C, 0x1E, 0x16, 0x1D, 0x2F, 0x59, 0x5B, 0x24, 0x59,
	0x2E, 0x08, 0x52, 0x11, 0x29, 0x18, 0x1E, 0x3F, 0x74, 0x15, 0x32, 0x18,
	0x11, 0x21, 0x16, 0x55, 0x45, 0x3F, 0x32, 0x03, 0x0C, 0x1A, 0x01, 0x04,
	0x1D, 0x58, 0x3B, 0x5B, 0x13, 0x2B, 0x34, 0x02, 0x18, 0x14, 0x1A, 0x2D,
	0x3D, 0x08, 0x05, 0x22, 0x38, 0x3C, 0x26, 0x35, 0x16, 0x13, 0x20, 0x1B,
	0x23, 0x18, 0x39, 0x2C, 0x1D, 0x2E, 0x2A, 0x56, 0x3E, 0x11, 0x38, 0x09,
	0x2E, 0x3A, 0x23, 0x28, 0x18, 0x02, 0x1A, 0x5A, 0x29, 0x1E, 0x1B, 0x28,
	0x27, 0x2E, 0x0A, 0x3B, 0x41, 0x26, 0x07, 0x07, 0x12, 0x39, 0x3A, 0x6D,
	0x2D, 0x00, 0x2D, 0x00, 0x07, 0x3E, 0x4E, 0x39, 0x00, 0x28, 0x5C, 0x00,
	0x1B, 0x0F, 0x15, 0x20, 0x18, 0x03, 0x59, 0x25, 0x0F, 0x37, 0x0A, 0x21,
	0x2E, 0x0B, 0x11, 0x00, 0x2D, 0x7B, 0x2A, 0x50, 0x58, 0x1A, 0x0B, 0x1C,
	0x3B, 0x14, 0x2E, 0x0E, 0x1F, 0x0A, 0x2A, 0x59, 0x10, 0x0D, 0x23, 0x08,
	0x0A, 0x2E, 0x19, 0x4A, 0x41, 0x1F, 0x01, 0x23, 0x2F, 0x18, 0x11, 0x24,
	0x02, 0x0D, 0x5F, 0x07, 0x36, 0x58, 0x19, 0x27, 0x08, 0x13, 0x1B, 0x30,
	0x5B, 0x3D, 0x7B, 0x36, 0x30, 0x36, 0x23, 0x14, 0x07, 0x38, 0x5E, 0x5C,
	0x24, 0x54, 0x25, 0x41, 0x39, 0x24, 0x47, 0x09, 0x2C, 0x28, 0x2E, 0x5B,
	0x0A, 0x56, 0x58, 0x2B, 0x23, 0x2F, 0x2A, 0x02, 0x6D, 0x25, 0x0F, 0x02,
	0x59, 0x2D, 0x0E, 0x05, 0x05, 0x0E, 0x38, 0x54, 0x27, 0x05, 0x09, 0x34,
	0x21, 0x2C, 0x3E, 0x22, 0x75, 0x5E, 0x13, 0x3D, 0x00, 0x75, 0x54, 0x03,
	0x02, 0x2F, 0x31, 0x24, 0x24, 0x3E, 0x3B, 0x0E, 0x06, 0x23, 0x03, 0x53,
	0x35, 0x23, 0x32, 0x3C, 0x1E, 0x0D, 0x20, 0x28, 0x1F, 0x18, 0x17, 0x5B,
	0x05, 0x17, 0x5E, 0x27, 0x08, 0x36, 0x3D, 0x3E, 0x72, 0x01, 0x04, 0x0C,
	0x03, 0x01, 0x16, 0x2C, 0x1E, 0x08, 0x0E, 0x35, 0x30, 0x21, 0x58, 0x1B,
	0x5F, 0x32, 0x22, 0x1B, 0x17, 0x22, 0x0D, 0x23, 0x08, 0x12, 0x35, 0x2C,
	0x36, 0x00, 0x2E, 0x47, 0x05, 0x38, 0x40, 0x2B, 0x0D, 0x22, 0x02, 0x11,
	0x1A, 0x2F, 0x2B, 0x0F, 0x2E, 0x2A, 0x5F, 0x29, 0x09, 0x25, 0x15, 0x1E,
	0x52, 0x3B, 0x23, 0x2F, 0x27, 0x4E, 0x14, 0x33, 0x7A, 0x55, 0x27, 0x5E,
	0x5C, 0x25, 0x5E, 0x2C, 0x14, 0x0A, 0x27, 0x38, 0x4A, 0x3F, 0x44, 0x2F,
	0x03, 0x55, 0x26, 0x58, 0x74, 0x01, 0x57, 0x5C, 0x2D, 0x35, 0x1E, 0x10,
	0x34, 0x1E, 0x3B, 0x0F, 0x20, 0x27, 0x28, 0x00, 0x0E, 0x36, 0x5F, 0x22,
	0x16, 0x1E, 0x06, 0x0B, 0x12, 0x7A, 0x0A, 0x51, 0x3F, 0x32, 0x0E, 0x0E,
	0x3B, 0x16, 0x5B, 0x0E, 0x27, 0x57, 0x3E, 0x06, 0x08, 0x0D, 0x26, 0x58,
	0x18, 0x3A, 0x1D, 0x15, 0x02, 0x1E, 0x69, 0x1D, 0x06, 0x5C, 0x02, 0x08,
	0x1E, 0x37, 0x41, 0x13, 0x01, 0x5D, 0x29, 0x05, 0x28, 0x20, 0x2E, 0x04,
	0x3C, 0x23, 0x2C, 0x14, 0x02, 0x05, 0x13, 0x17, 0x1A, 0x31, 0x3D, 0x1C,
	0x30, 0x2F, 0x15, 0x2D, 0x0D, 0x14, 0x47, 0x34, 0x0D, 0x5D, 0x75, 0x35,
	0x35, 0x36, 0x1F, 0x34, 0x5E, 0x23, 0x3C, 0x5B, 0x1B, 0x0E, 0x51, 0x22,
	0x5B, 0x18, 0x0D, 0x15, 0x04, 0x40, 0x16, 0x55, 0x04, 0x21, 0x0A, 0x3A,
	0x39, 0x28, 0x09, 0x0A, 0x29, 0x09, 0x35, 0x08, 0x3C, 0x11, 0x21, 0x4A,
	0x0F, 0x18, 0x10, 0x28, 0x25, 0x5E, 0x1F, 0x18, 0x39, 0x30, 0x57, 0x21,
	0x0A, 0x1A, 0x0B, 0x26, 0x27, 0x31, 0x28, 0x20, 0x41, 0x5D, 0x04, 0x43,
	0x04, 0x00, 0x2E, 0x14, 0x15, 0x57, 0x5D, 0x38, 0x21, 0x07, 0x53, 0x07,
	0x5A, 0x77, 0x22, 0x50, 0x05, 0x04, 0x38, 0x2F, 0x1B, 0x38, 0x02, 0x2D,
	0x3A, 0x11, 0x21, 0x27, 0x06, 0x3F, 0x13, 0x1B, 0x0A, 0x13, 0x08, 0x52,
	0x16, 0x08, 0x34, 0x28, 0x0C, 0x16, 0x33, 0x69, 0x1D, 0x37, 0x5C, 0x22,
	0x14, 0x47, 0x14, 0x3C, 0x26, 0x73, 0x14, 0x2A, 0x00, 0x0C, 0x17, 0x3D,
	0x32, 0x1F, 0x07, 0x32, 0x04, 0x1B, 0x2B, 0x13, 0x2E, 0x05, 0x28, 0x2F,
	0x2F, 0x03, 0x21, 0x50, 0x58, 0x3D, 0x13, 0x09, 0x33, 0x19, 0x44, 0x03,
	0x0D, 0x13, 0x56, 0x53, 0x71, 0x26, 0x55, 0x0B, 0x5F, 0x37, 0x3F, 0x35,
	0x2C, 0x21, 0x32, 0x34, 0x1B, 0x21, 0x0A, 0x01, 0x03, 0x3B, 0x1C, 0x32,
	0x29, 0x2D, 0x4E, 0x06, 0x07, 0x0B, 0x0A, 0x00, 0x00, 0x2F, 0x00, 0x5B,
	0x2B, 0x0B, 0x05, 0x7B, 0x43, 0x24, 0x3C, 0x04, 0x10, 0x59, 0x31, 0x04,
	0x44, 0x31, 0x35, 0x0A, 0x39, 0x1C, 0x18, 0x25, 0x0A, 0x59, 0x3D, 0x70,
	0x08, 0x25, 0x5D, 0x2D, 0x2D, 0x5F, 0x12, 0x0A, 0x5D, 0x77, 0x55, 0x09,
	0x09, 0x12, 0x2F, 0x35, 0x30, 0x18, 0x20, 0x1B, 0x03, 0x30, 0x06, 0x27,
	0x10, 0x20, 0x18, 0x1B, 0x13, 0x2C, 0x5B, 0x39, 0x3C, 0x07, 0x73, 0x23,
	0x51, 0x21, 0x53, 0x74, 0x5D, 0x15, 0x5D, 0x00, 0x06, 0x59, 0x13, 0x14,
	0x40, 0x3A, 0x1D, 0x02, 0x06, 0x0A, 0x0B, 0x05, 0x20, 0x1A, 0x21, 0x17,
	0x36, 0x58, 0x08, 0x0A, 0x1B, 0x3B, 0x0E, 0x1A, 0x2A, 0x34, 0x1E, 0x2E,
	0x29, 0x07, 0x36, 0x1F, 0x2B, 0x36, 0x5C, 0x17, 0x47, 0x2C, 0x3B, 0x3F,
	0x10, 0x15, 0x39, 0x2F, 0x0C, 0x1B, 0x14, 0x10, 0x5E, 0x0F, 0x31, 0x02,
	0x51, 0x39, 0x0A, 0x32, 0x27, 0x04, 0x5A, 0x2C, 0x2D, 0x04, 0x20, 0x14,
	0x21, 0x34, 0x09, 0x51, 0x39, 0x0E, 0x32, 0x35, 0x57, 0x27, 0x2A, 0x35,
	0x1F, 0x14, 0x16, 0x24, 0x0F, 0x2A, 0x0B, 0x18, 0x27, 0x0E, 0x0A, 0x2D,
	0x5C, 0x5F, 0x08, 0x0A, 0x12, 0x26, 0x2C, 0x28, 0x19, 0x3B, 0x1A, 0x1D,
	0x76, 0x21, 0x08, 0x02, 0x29, 0x04, 0x0E, 0x08, 0x1F, 0x59, 0x2F, 0x5F,
	0x26, 0x3F, 0x02, 0x29, 0x07, 0x14, 0x16, 0x24, 0x05, 0x5C, 0x59, 0x41,
	0x2C, 0x3B, 0x3F, 0x17, 0x03, 0x5A, 0x0B, 0x00, 0x04, 0x39, 0x5C, 0x23,
	0x3D, 0x4E, 0x3F, 0x2E, 0x16, 0x0E, 0x29, 0x2D, 0x05, 0x18, 0x35, 0x27,
	0x18, 0x5B, 0x71, 0x1D, 0x0E, 0x59, 0x58, 0x73, 0x5F, 0x2C, 0x19, 0x0D,
	0x70, 0x25, 0x12, 0x2A, 0x25, 0x24, 0x2F, 0x37, 0x19, 0x5B, 0x05, 0x5D,
	0x1B, 0x2B, 0x23, 0x2E, 0x16, 0x50, 0x3D, 0x53, 0x2E, 0x5D, 0x0F, 0x01,
	0x07, 0x6D, 0x36, 0x0C, 0x00, 0x2D, 0x08, 0x2D, 0x2C, 0x16, 0x58, 0x27,
	0x3C, 0x1B, 0x02, 0x28, 0x04, 0x1A, 0x11, 0x34, 0x0C, 0x04, 0x20, 0x38,
	0x0A, 0x5D, 0x38, 0x55, 0x25, 0x3F, 0x59, 0x7A, 0x0B, 0x06, 0x5D, 0x53,
	0x21, 0x3D, 0x30, 0x0C, 0x1E, 0x03, 0x1B, 0x00, 0x2D, 0x2F, 0x20, 0x29,
	0x53, 0x5C, 0x40, 0x29, 0x1A, 0x55, 0x3E, 0x40, 0x21, 0x14, 0x23, 0x34,
	0x39, 0x26, 0x5C, 0x4E, 0x21, 0x1D, 0x32, 0x2D, 0x35, 0x18, 0x26, 0x6D,
	0x24, 0x04, 0x19, 0x0C, 0x32, 0x16, 0x17, 0x5A, 0x40, 0x17, 0x2D, 0x2F,
	0x2C, 0x2F, 0x2D, 0x27, 0x04, 0x41, 0x1D, 0x74, 0x3A, 0x2F, 0x03, 0x3E,
	0x0B, 0x1A, 0x2F, 0x01, 0x29, 0x20, 0x07, 0x03, 0x2A, 0x27, 0x35, 0x1A,
	0x2E, 0x1B, 0x18, 0x18, 0x43, 0x51, 0x3B, 0x06, 0x33, 0x22, 0x2E, 0x1A,
	0x2A, 0x70, 0x02, 0x0C, 0x3E, 0x2C, 0x75, 0x3A, 0x50, 0x37, 0x29, 0x18,
	0x1C, 0x56, 0x21, 0x5E, 0x15, 0x0B, 0x1B, 0x21, 0x24, 0x32, 0x1F, 0x18,
	0x37, 0x01, 0x3B, 0x3B, 0x2F, 0x39, 0x23, 0x18, 0x28, 0x14, 0x3B, 0x32,
	0x13, 0x15, 0x0D, 0x1E, 0x1C, 0x3B, 0x3B, 0x3B, 0x5E, 0x01, 0x71, 0x05,
	0x4E, 0x39, 0x1E, 0x70, 0x27, 0x35, 0x08, 0x07, 0x15, 0x03, 0x36, 0x02,
	0x04, 0x73, 0x25, 0x2A, 0x05, 0x3D, 0x0D, 0x3A, 0x2E, 0x0D, 0x32, 0x17,
	0x0B, 0x2A, 0x38, 0x1E, 0x36, 0x1F, 0x11, 0x20, 0x3D, 0x30, 0x00, 0x26,
	0x36, 0x18, 0x24, 0x54, 0x31, 0x56, 0x32, 0x04, 0x5D, 0x16, 0x2C, 0x2E,
	0x20, 0x07, 0x2D, 0x0A, 0x1D, 0x74, 0x3D, 0x22, 0x2B, 0x32, 0x0B, 0x0D,
	0x20, 0x5D, 0x1D, 0x7A, 0x20, 0x28, 0x5D, 0x58, 0x16, 0x3E, 0x32, 0x28,
	0x21, 0x71, 0x16, 0x55, 0x34, 0x52, 0x0C, 0x29, 0x55, 0x3A, 0x23, 0x6D,
	0x3E, 0x2E, 0x26, 0x05, 0x0F, 0x1D, 0x27, 0x36, 0x0C, 0x33, 0x0D, 0x2E,
	0x01, 0x53, 0x0C, 0x25, 0x39, 0x01, 0x0E, 0x37, 0x2B, 0x00, 0x41, 0x13,
	0x12, 0x01, 0x16, 0x26, 0x40, 0x17, 0x00, 0x16, 0x0F, 0x39, 0x2B, 0x0B,
	0x4E, 0x41, 0x0D, 0x73, 0x38, 0x53, 0x58, 0x44, 0x6D, 0x02, 0x0C, 0x5A,
	0x44, 0x2D, 0x08, 0x11, 0x41, 0x33, 0x26, 0x1E, 0x57, 0x5B, 0x44, 0x0F,
	0x5D, 0x0B, 0x56, 0x1B, 0x34, 0x3C, 0x57, 0x26, 0x3A, 0x12, 0x23, 0x2B,
	0x22, 0x05, 0x74, 0x54, 0x07, 0x19, 0x5D, 0x28, 0x05, 0x2C, 0x5B, 0x06,
	0x17, 0x3E, 0x2C, 0x5C, 0x02, 0x31, 0x1D, 0x19, 0x26, 0x3A, 0x25, 0x0E,
	0x23, 0x2C, 0x2C, 0x09, 0x0F, 0x0C, 0x1D, 0x28, 0x2A, 0x23, 0x0F, 0x1C,
	0x07, 0x25, 0x0E, 0x23, 0x41, 0x39, 0x72, 0x06, 0x18, 0x28, 0x53, 0x0D,
	0x07, 0x22, 0x56, 0x22, 0x11, 0x3F, 0x16, 0x1D, 0x3B, 0x38, 0x1D, 0x09,
	0x23, 0x5E, 0x13, 0x0A, 0x39, 0x1B, 0x25, 0x17, 0x2B, 0x22, 0x09, 0x20,
	0x29, 0x25, 0x0B, 0x27, 0x5D, 0x0E, 0x22, 0x2F, 0x39, 0x23, 0x32, 0x38,
	0x22, 0x1B, 0x19, 0x38, 0x1E, 0x0D, 0x0F, 0x52, 0x76, 0x5E, 0x54, 0x01,
	0x5C, 0x2C, 0x00, 0x0E, 0x2A, 0x00, 0x32, 0x09, 0x0A, 0x37, 0x08, 0x3B,
	0x1A, 0x2C, 0x28, 0x5E, 0x35, 0x0F, 0x33, 0x3D, 0x20, 0x04, 0x39, 0x07,
	0x18, 0x2F, 0x03, 0x2B, 0x39, 0x45, 0x3B, 0x2E, 0x39, 0x18, 0x3E, 0x03,
	0x72, 0x5E, 0x06, 0x01, 0x3D, 0x03, 0x2E, 0x02, 0x26, 0x1A, 0x06, 0x3E,
	0x31, 0x19, 0x53, 0x73, 0x5E, 0x37, 0x1E, 0x12, 0x0F, 0x1B, 0x37, 0x0B,
	0x21, 0x09, 0x58, 0x59, 0x05, 0x44, 0x04, 0x22, 0x55, 0x5A, 0x2C, 0x30,
	0x2D, 0x32, 0x1D, 0x58, 0x31, 0x5B, 0x24, 0x0D, 0x1D, 0x0E, 0x1E, 0x58,
	0x39, 0x24, 0x2D, 0x20, 0x09, 0x25, 0x3E, 0x28, 0x39, 0x06, 0x01, 0x29,
	0x23, 0x18, 0x58, 0x34, 0x33, 0x11, 0x5D, 0x57, 0x19, 0x0D, 0x0F, 0x58,
	0x30, 0x2C, 0x39, 0x09, 0x20, 0x0E, 0x29, 0x38, 0x25, 0x0F, 0x0A, 0x3C,
	0x40, 0x3B, 0x29, 0x16, 0x1C, 0x28, 0x73, 0x23, 0x30, 0x41, 0x5F, 0x6D,
	0x1E, 0x4A, 0x0A, 0x09, 0x12, 0x08, 0x14, 0x1A, 0x5E, 0x76, 0x2A, 0x09,
	0x1D, 0x21, 0x76, 0x38, 0x25, 0x1B, 0x21, 0x74, 0x0A, 0x15, 0x04, 0x22,
	0x73, 0x1A, 0x31, 0x0B, 0x05, 0x34, 0x24, 0x51, 0x18, 0x2F, 0x1A, 0x58,
	0x05, 0x41, 0x3A, 0x7A, 0x24, 0x24, 0x0F, 0x18, 0x32, 0x00, 0x24, 0x2A,
	0x44, 0x76, 0x29, 0x26, 0x01, 0x0C, 0x37, 0x3C, 0x4E, 0x24, 0x0E, 0x32,
	0x2F, 0x56, 0x04, 0x52, 0x12, 0x29, 0x13, 0x28, 0x2D, 0x21, 0x5E, 0x56,
	0x03, 0x39, 0x74, 0x1C, 0x30, 0x45, 0x06, 0x10, 0x07, 0x55, 0x0D, 0x3B,
	0x2F, 0x0E, 0x58, 0x29, 0x13, 0x13, 0x05, 0x30, 0x28, 0x23, 0x32, 0x26,
	0x1B, 0x38, 0x2F, 0x10, 0x47, 0x32, 0x03, 0x5F, 0x00, 0x14, 0x31, 0x14,
	0x3B, 0x3A, 0x1E, 0x53, 0x08, 0x20, 0x2D, 0x1A, 0x26, 0x3A, 0x2E, 0x75,
	0x1C, 0x4E, 0x38, 0x58, 0x33, 0x02, 0x0C, 0x25, 0x28, 0x37, 0x0A, 0x58,
	0x56, 0x3F, 0x37, 0x1C, 0x38, 0x5A, 0x21, 0x75, 0x2A, 0x18, 0x5F, 0x3C,
	0x71, 0x19, 0x13, 0x3C, 0x29, 0x32, 0x2F, 0x39, 0x1A, 0x32, 0x1A, 0x36,
	0x53, 0x59, 0x25, 0x7B, 0x14, 0x31, 0x57, 0x13, 0x35, 0x5C, 0x35, 0x36,
	0x22, 0x37, 0x2B, 0x4A, 0x02, 0x21, 0x0B, 0x0F, 0x37, 0x1F, 0x31, 0x72,
	0x22, 0x3B, 0x24, 0x07, 0x1A, 0x34, 0x24, 0x1B, 0x26, 0x03, 0x3D, 0x16,
	0x0D, 0x1A, 0x0B, 0x23, 0x26, 0x1F, 0x32, 0x0F, 0x08, 0x30, 0x26, 0x24,
	0x1A, 0x2F, 0x56, 0x39, 0x1A, 0x23, 0x59, 0x26, 0x23, 0x3B, 0x2E, 0x0E,
	0x06, 0x3E, 0x19, 0x30, 0x0B, 0x32, 0x59, 0x27, 0x29, 0x27, 0x2A, 0x06,
	0x3E, 0x36, 0x29, 0x0C, 0x1B, 0x5D, 0x75, 0x0F, 0x57, 0x06, 0x59, 0x2A,
	0x3D, 0x58, 0x17, 0x5A, 0x0C, 0x2E, 0x36, 0x57, 0x21, 0x7A, 0x07, 0x56,
	0x3C, 0x0D, 0x6D, 0x47, 0x2B, 0x28, 0x0D, 0x27, 0x23, 0x23, 0x07, 0x21,
	0x0A, 0x1F, 0x00, 0x00, 0x58, 0x35, 0x16, 0x57, 0x18, 0x39, 0x37, 0x04,
	0x06, 0x59, 0x1D, 0x77, 0x55, 0x59, 0x26, 0x26, 0x0A, 0x58, 0x28, 0x0D,
	0x32, 0x25, 0x35, 0x0E, 0x3C, 0x2C, 0x01, 0x5E, 0x52, 0x22, 0x05, 0x29,
	0x25, 0x03, 0x05, 0x3E, 0x0D, 0x21, 0x37, 0x34, 0x32, 0x2B, 0x3A, 0x4E,
	0x2D, 0x2D, 0x10, 0x34, 0x05, 0x2D, 0x0C, 0x13, 0x28, 0x14, 0x26, 0x0E,
	0x1B, 0x14, 0x57, 0x29, 0x1E, 0x29, 0x59, 0x14, 0x09, 0x1A, 0x3A, 0x0D,
	0x1B, 0x27, 0x20, 0x1A, 0x0F, 0x2B, 0x37, 0x19, 0x75, 0x54, 0x09, 0x45,
	0x5C, 0x09, 0x3B, 0x32, 0x36, 0x5C, 0x01, 0x26, 0x00, 0x08, 0x2E, 0x0D,
	0x06, 0x29, 0x08, 0x5D, 0x01, 0x03, 0x0E, 0x28, 0x2D, 0x72, 0x08, 0x05,
	0x16, 0x28, 0x24, 0x3A, 0x22, 0x0F, 0x2A, 0x0A, 0x2E, 0x29, 0x5A, 0x28,
	0x73, 0x26, 0x26, 0x3E, 0x04, 0x20, 0x5D, 0x52, 0x28, 0x0A, 0x3A, 0x3D,
	0x53, 0x3C, 0x05, 0x3B, 0x2B, 0x58, 0x19, 0x3B, 0x04, 0x0F, 0x0A, 0x5E,
	0x32, 0x24, 0x04, 0x0D, 0x18, 0x0F, 0x14, 0x5A, 0x32, 0x56, 0x12, 0x27,
	0x5D, 0x34, 0x21, 0x02, 0x0C, 0x5E, 0x07, 0x28, 0x0D, 0x28, 0x5F, 0x03,
	0x1D, 0x52, 0x2D, 0x0B, 0x4A, 0x01, 0x53, 0x03, 0x3A, 0x03, 0x37, 0x1C,
	0x0F, 0x0F, 0x14, 0x3A, 0x03, 0x21, 0x58, 0x02, 0x03, 0x04, 0x1B, 0x27,
	0x02, 0x0A, 0x03, 0x3B, 0x59, 0x14, 0x0D, 0x2F, 0x2D, 0x15, 0x29, 0x41,
	0x52, 0x76, 0x59, 0x4A, 0x3E, 0x18, 0x34, 0x15, 0x12, 0x22, 0x1C, 0x36,
	0x3D, 0x56, 0x03, 0x58, 0x0D, 0x15, 0x11, 0x18, 0x21, 0x15, 0x3A, 0x16,
	0x20, 0x0D, 0x2E, 0x3C, 0x03, 0x3B, 0x1A, 0x2A, 0x3B, 0x04, 0x3D, 0x39,
	0x71, 0x58, 0x0A, 0x2A, 0x06, 0x17, 0x2D, 0x29, 0x38, 0x1D, 0x1B, 0x5C,
	0x0E, 0x1B, 0x39, 0x35, 0x24, 0x26, 0x57, 0x1F, 0x03, 0x28, 0x24, 0x1F,
	0x0E, 0x11, 0x08, 0x1B, 0x03, 0x5E, 0x28, 0x18, 0x06, 0x20, 0x3C, 0x76,
	0x2E, 0x0B, 0x34, 0x1D, 0x24, 0x58, 0x31, 0x20, 0x3E, 0x2E, 0x43, 0x59,
	0x29, 0x24, 0x31, 0x3C, 0x0D, 0x3D, 0x12, 0x3B, 0x3A, 0x32, 0x3E, 0x20,
	0x13, 0x29, 0x36, 0x1D, 0x0F, 0x03, 0x2E, 0x35, 0x17, 0x3B, 0x25, 0x47,
	0x1B, 0x2D, 0x0F, 0x76, 0x38, 0x0A, 0x3A, 0x44, 0x28, 0x59, 0x02, 0x3E,
	0x06, 0x28, 0x59, 0x30, 0x34, 0x02, 0x34, 0x14, 0x0A, 0x34, 0x02, 0x0C,
	0x1D, 0x06, 0x39, 0x3D, 0x00, 0x1E, 0x33, 0x22, 0x3A, 0x0D, 0x2B, 0x13,
	0x22, 0x58, 0x33, 0x38, 0x33, 0x03, 0x28, 0x16, 0x2F, 0x59, 0x5D, 0x2A,
	0x3B, 0x0B, 0x17, 0x59, 0x27, 0x28, 0x25, 0x28, 0x00, 0x05, 0x21, 0x3F,
	0x00, 0x2C, 0x0D, 0x0C, 0x3A, 0x36, 0x3B, 0x2A, 0x71, 0x0A, 0x27, 0x1D,
	0x5D, 0x77, 0x16, 0x22, 0x18, 0x1A, 0x09, 0x1F, 0x15, 0x09, 0x3B, 0x17,
	0x0E, 0x30, 0x16, 0x3A, 0x2B, 0x59, 0x08, 0x0D, 0x2A, 0x29, 0x2F, 0x05,
	0x1D, 0x5C, 0x69, 0x06, 0x31, 0x0C, 0x00, 0x2D, 0x2E, 0x0A, 0x5A, 0x02,
	0x21, 0x2D, 0x0B, 0x29, 0x22, 0x07, 0x38, 0x34, 0x0C, 0x40, 0x15, 0x5B,
	0x51, 0x1D, 0x09, 0x1B, 0x1A, 0x26, 0x45, 0x05, 0x0F, 0x0A, 0x52, 0x41,
	0x25, 0x3A, 0x19, 0x15, 0x2C, 0x1F, 0x01, 0x15, 0x11, 0x2D, 0x59, 0x08,
	0x1C, 0x2D, 0x16, 0x25, 0x29, 0x5B, 0x34, 0x1E, 0x27, 0x37, 0x0E, 0x39,
	0x25, 0x2E, 0x28, 0x20, 0x15, 0x38, 0x00, 0x33, 0x2E, 0x07, 0x0D, 0x13,
	0x18, 0x2D, 0x32, 0x25, 0x0A, 0x26, 0x29, 0x4A, 0x5B, 0x2E, 0x71, 0x5D,
	0x12, 0x08, 0x5F, 0x00, 0x0D, 0x37, 0x04, 0x18, 0x37, 0x03, 0x08, 0x16,
	0x0E, 0x32, 0x2F, 0x24, 0x0B, 0x03, 0x01, 0x1F, 0x32, 0x5B, 0x32, 0x26,
	0x03, 0x05, 0x26, 0x28, 0x7B, 0x27, 0x23, 0x36, 0x2F, 0x05, 0x3D, 0x53,
	0x2D, 0x40, 0x76, 0x34, 0x36, 0x24, 0x3B, 0x28, 0x55, 0x0C, 0x02, 0x59,
	0x2E, 0x1B, 0x50, 0x3F, 0x3C, 0x21, 0x1D, 0x06, 0x08, 0x39, 0x2B, 0x43,
	0x22, 0x1D, 0x3B, 0x3B, 0x04, 0x50, 0x5E, 0x2D, 0x21, 0x16, 0x07, 0x06,
	0x00, 0x01, 0x38, 0x0D, 0x29, 0x40, 0x38, 0x24, 0x09, 0x05, 0x20, 0x34,
	0x15, 0x05, 0x05, 0x1D, 0x2F, 0x2E, 0x13, 0x03, 0x2D, 0x71, 0x35, 0x53,
	0x2A, 0x1F, 0x37, 0x1B, 0x0C, 0x39, 0x1C, 0x21, 0x29, 0x0E, 0x59, 0x2F,
	0x08, 0x06, 0x04, 0x09, 0x12, 0x72, 0x2E, 0x1B, 0x28, 0x52, 0x35, 0x2D,
	0x51, 0x06, 0x00, 0x72, 0x25, 0x31, 0x25, 0x23, 0x1B, 0x28, 0x32, 0x5A,
	0x19, 0x23, 0x3F, 0x37, 0x1A, 0x20, 0x11, 0x59, 0x0D, 0x2F, 0x20, 0x76,
	0x2E, 0x0F, 0x3A, 0x32, 0x08, 0x20, 0x0B, 0x59, 0x2C, 0x72, 0x0B, 0x08,
	0x02, 0x24, 0x7A, 0x00, 0x00, 0x17, 0x06, 0x09, 0x0A, 0x54, 0x1E, 0x1A,
	0x12, 0x05, 0x15, 0x29, 0x23, 0x25, 0x2F, 0x56, 0x36, 0x0F, 0x21, 0x54,
	0x0E, 0x1F, 0x52, 0x00, 0x0F, 0x29, 0x0D, 0x05, 0x0D, 0x5E, 0x33, 0x1D,
	0x3C, 0x30, 0x1C, 0x2F, 0x29, 0x3C, 0x26, 0x2B, 0x2B, 0x5C, 0x1C, 0x12,
	0x27, 0x53, 0x38, 0x5F, 0x69, 0x2D, 0x33, 0x1F, 0x07, 0x34, 0x16, 0x36,
	0x05, 0x44, 0x20, 0x2B, 0x55, 0x1C, 0x3B, 0x0F, 0x5E, 0x08, 0x1D, 0x21,
	0x36, 0x5D, 0x04, 0x28, 0x5C, 0x13, 0x5D, 0x04, 0x25, 0x12, 0x0E, 0x5E,
	0x57, 0x1D, 0x1B, 0x07, 0x2B, 0x2F, 0x21, 0x27, 0x71, 0x5E, 0x2E, 0x1C,
	0x53, 0x2B, 0x2A, 0x2B, 0x5D, 0x00, 0x0D, 0x25, 0x20, 0x03, 0x0A, 0x25,
	0x08, 0x16, 0x45, 0x24, 0x74, 0x0B, 0x23, 0x1B, 0x2E, 0x20, 0x04, 0x36,
	0x3E, 0x13, 0x16, 0x09, 0x54, 0x1C, 0x3F, 0x27, 0x35, 0x56, 0x5E, 0x58,
	0x72, 0x2D, 0x59, 0x5E, 0x05, 0x6D, 0x2F, 0x2A, 0x45, 0x39, 0x37, 0x5B,
	0x53, 0x5D, 0x39, 0x69, 0x23, 0x56, 0x1F, 0x01, 0x26, 0x15, 0x05, 0x24,
	0x08, 0x32, 0x5F, 0x06, 0x16, 0x1F, 0x00, 0x19, 0x51, 0x2F, 0x23, 0x6D,
	0x28, 0x10, 0x07, 0x5F, 0x34, 0x47, 0x55, 0x0B, 0x07, 0x09, 0x2F, 0x23,
	0x27, 0x3F, 0x15, 0x2E, 0x16, 0x2C, 0x11, 0x31, 0x1B, 0x02, 0x34, 0x27,
	0x7B, 0x07, 0x0A, 0x37, 0x12, 0x08, 0x0D, 0x3B, 0x14, 0x2F, 0x75, 0x3E,
	0x20, 0x2F, 0x1F, 0x2B, 0x1D, 0x51, 0x1E, 0x20, 0x37, 0x21, 0x0D, 0x1D,
	0x1F, 0x6D, 0x1B, 0x12, 0x1B, 0x3B, 0x70, 0x03, 0x03, 0x01, 0x3F, 0x7B,
	0x07, 0x04, 0x5B, 0x19, 0x25, 0x22, 0x3B, 0x3F, 0x28, 0x10, 0x34, 0x02,
	0x1A, 0x21, 0x05, 0x05, 0x54, 0x24, 0x18, 0x10, 0x3D, 0x2F, 0x1C, 0x53,
	0x77, 0x01, 0x29, 0x2B, 0x3E, 0x24, 0x36, 0x53, 0x5C, 0x18, 0x13, 0x54,
	0x24, 0x3E, 0x23, 0x08, 0x16, 0x2F, 0x0A, 0x23, 0x24, 0x28, 0x2A, 0x1A,
	0x11, 0x01, 0x0A, 0x0B, 0x26, 0x0F, 0x0A, 0x03, 0x03, 0x5E, 0x07, 0x35,
	0x47, 0x02, 0x2C, 0x0E, 0x21, 0x1D, 0x32, 0x02, 0x12, 0x70, 0x3B, 0x32,
	0x08, 0x2D, 0x16, 0x18, 0x07, 0x19, 0x03, 0x2C, 0x09, 0x57, 0x5D, 0x31,
	0x32, 0x0B, 0x2F, 0x19, 0x20, 0x27, 0x5D, 0x0E, 0x5A, 0x02, 0x0E, 0x2D,
	0x10, 0x2F, 0x38, 0x03, 0x3A, 0x26, 0x08, 0x59, 0x1B, 0x2F, 0x19, 0x0A,
	0x5F, 0x0B, 0x1D, 0x2F, 0x2F, 0x3E, 0x32, 0x47, 0x03, 0x14, 0x0F, 0x37,
	0x2E, 0x10, 0x2A, 0x39, 0x70, 0x00, 0x53, 0x3B, 0x3F, 0x11, 0x43, 0x09,
	0x03, 0x5B, 0x23, 0x00, 0x54, 0x2F, 0x25, 0x76, 0x19, 0x06, 0x5D, 0x5C,
	0x05, 0x01, 0x02, 0x21, 0x59, 0x05, 0x0B, 0x58, 0x0A, 0x0C, 0x0F, 0x02,
	0x18, 0x0C, 0x00, 0x01, 0x23, 0x24, 0x02, 0x3D, 0x01, 0x47, 0x51, 0x20,
	0x58, 0x1B, 0x5A, 0x4E, 0x1E, 0x40, 0x73, 0x28, 0x13, 0x1C, 0x20, 0x3B,
	0x0B, 0x04, 0x0B, 0x22, 0x2E, 0x2D, 0x2E, 0x5B, 0x1B, 0x0B, 0x02, 0x24,
	0x3A, 0x38, 0x3A, 0x3C, 0x50, 0x5D, 0x5E, 0x2B, 0x1E, 0x06, 0x20, 0x06,
	0x24, 0x5E, 0x14, 0x2D, 0x0F, 0x76, 0x3D, 0x3B, 0x16, 0x3C, 0x04, 0x2D,
	0x27, 0x3F, 0x52, 0x2B, 0x3C, 0x56, 0x04, 0x53, 0x20, 0x29, 0x54, 0x16,
	0x2F, 0x00, 0x24, 0x11, 0x41, 0x25, 0x0E, 0x08, 0x29, 0x08, 0x33, 0x10,
	0x23, 0x2D, 0x01, 0x2F, 0x69, 0x23, 0x35, 0x2A, 0x0D, 0x0C, 0x2D, 0x04,
	0x2F, 0x02, 0x0D, 0x54, 0x08, 0x0D, 0x58, 0x0A, 0x06, 0x53, 0x45, 0x3D,
	0x00, 0x03, 0x13, 0x37, 0x2F, 0x1A, 0x14, 0x56, 0x06, 0x02, 0x73, 0x3C,
	0x13, 0x1F, 0x3F, 0x25, 0x16, 0x0E, 0x5B, 0x02, 0x70, 0x03, 0x54, 0x39,
	0x00, 0x23, 0x34, 0x32, 0x0B, 0x3E, 0x07, 0x2D, 0x30, 0x41, 0x1C, 0x2C,
	0x3E, 0x14, 0x00, 0x1B, 0x0E, 0x3B, 0x1B, 0x08, 0x3B, 0x37, 0x14, 0x56,
	0x0C, 0x2D, 0x7B, 0x1B, 0x1B, 0x17, 0x0A, 0x15, 0x3A, 0x04, 0x08, 0x53,
	0x1A, 0x3A, 0x2B, 0x3D, 0x13, 0x72, 0x21, 0x37, 0x1B, 0x59, 0x27, 0x5B,
	0x59, 0x57, 0x11, 0x03, 0x39, 0x0D, 0x0F, 0x07, 0x25, 0x21, 0x10, 0x04,
	0x3B, 0x7B, 0x27, 0x2E, 0x56, 0x2D, 0x30, 0x25, 0x33, 0x3D, 0x04, 0x15,
	0x43, 0x36, 0x5B, 0x0F, 0x25, 0x3F, 0x06, 0x3D, 0x0D, 0x0C, 0x3E, 0x26,
	0x0B, 0x00, 0x73, 0x3F, 0x12, 0x1B, 0x03, 0x18, 0x27, 0x56, 0x14, 0x32,
	0x06, 0x36, 0x27, 0x2B, 0x19, 0x25, 0x0A, 0x57, 0x3C, 0x22, 0x10, 0x29,
	0x26, 0x09, 0x3C, 0x29, 0x5D, 0x2D, 0x2D, 0x1B, 0x17, 0x55, 0x16, 0x23,
	0x27, 0x03, 0x08, 0x55, 0x09, 0x05, 0x73, 0x0D, 0x09, 0x5E, 0x18, 0x00,
	0x1B, 0x4A, 0x09, 0x0D, 0x21, 0x26, 0x25, 0x04, 0x21, 0x70, 0x26, 0x38,
	0x58, 0x3C, 0x04, 0x09, 0x38, 0x2B, 0x0D, 0x18, 0x3C, 0x36, 0x1B, 0x05,
	0x7B, 0x04, 0x57, 0x1A, 0x2C, 0x0C, 0x0D, 0x0B, 0x59, 0x58, 0x15, 0x3C,
	0x1B, 0x3C, 0x33, 0x13, 0x3D, 0x02, 0x1C, 0x3F, 0x2A, 0x5B, 0x39, 0x3C,
	0x18, 0x20, 0x24, 0x06, 0x5E, 0x23, 0x27, 0x25, 0x13, 0x03, 0x07, 0x32,
	0x5A, 0x02, 0x16, 0x5E, 0x0E, 0x34, 0x0B, 0x1B, 0x0C, 0x0F, 0x1D, 0x23,
	0x38, 0x5D, 0x03, 0x24, 0x20, 0x09, 0x1B, 0x2B, 0x3B, 0x00, 0x5A, 0x2E,
	0x69, 0x03, 0x56, 0x0D, 0x2E, 0x36, 0x04, 0x50, 0x2D, 0x06, 0x0F, 0x5E,
	0x57, 0x09, 0x26, 0x1A, 0x02, 0x57, 0x22, 0x1E, 0x2C, 0x5A, 0x37, 0x20,
	0x12, 0x0A, 0x3B, 0x23, 0x06, 0x25, 0x12, 0x03, 0x2C, 0x0A, 0x28, 0x21,
	0x07, 0x29, 0x5D, 0x3C, 0x2A, 0x1C, 0x29, 0x08, 0x00, 0x76, 0x2D, 0x2F,
	0x22, 0x32, 0x15, 0x15, 0x11, 0x36, 0x23, 0x11, 0x16, 0x18, 0x16, 0x5E,
	0x16, 0x08, 0x4E, 0x41, 0x03, 0x32, 0x3F, 0x56, 0x23, 0x0F, 0x76, 0x59,
	0x22, 0x2B, 0x32, 0x1B, 0x21, 0x17, 0x36, 0x39, 0x23, 0x20, 0x2B, 0x28,
	0x44, 0x1B, 0x3C, 0x59, 0x0A, 0x32, 0x72, 0x08, 0x50, 0x14, 0x05, 0x15,
	0x06, 0x53, 0x29, 0x3F, 0x73, 0x38, 0x06, 0x36, 0x5F, 0x26, 0x39, 0x4A,
	0x3B, 0x3B, 0x30, 0x19, 0x35, 0x3C, 0x2C, 0x14, 0x09, 0x59, 0x5F, 0x02,
	0x3B, 0x3F, 0x0C, 0x25, 0x20, 0x75, 0x05, 0x50, 0x45, 0x09, 0x32, 0x54,
	0x0F, 0x0B, 0x28, 0x18, 0x06, 0x56, 0x01, 0x24, 0x29, 0x26, 0x13, 0x00,
	0x2F, 0x7B, 0x1D, 0x08, 0x0D, 0x21, 0x04, 0x39, 0x0B, 0x25, 0x2F, 0x2E,
	0x47, 0x37, 0x2D, 0x1C, 0x2A, 0x1B, 0x06, 0x1D, 0x3A, 0x31, 0x1B, 0x16,
	0x2A, 0x08, 0x12, 0x14, 0x57, 0x38, 0x21, 0x6D, 0x5E, 0x28, 0x0C, 0x2F,
	0x06, 0x2B, 0x08, 0x25, 0x0C, 0x21, 0x36, 0x05, 0x2F, 0x00, 0x0C, 0x0D,
	0x28, 0x00, 0x5E, 0x2C, 0x36, 0x34, 0x01, 0x1E, 0x0C, 0x23, 0x09, 0x56,
	0x00, 0x32, 0x3F, 0x0B, 0x19, 0x11, 0x30, 0x5C, 0x2F, 0x1E, 0x31, 0x37,
	0x35, 0x55, 0x1C, 0x3D, 0x05, 0x2E, 0x52, 0x17, 0x5C, 0x38, 0x5C, 0x59,
	0x58, 0x25, 0x75, 0x5E, 0x3B, 0x25, 0x38, 0x2D, 0x0B, 0x11, 0x3C, 0x2E,
	0x14, 0x3C, 0x07, 0x58, 0x26, 0x0A, 0x00, 0x06, 0x2B, 0x27, 0x72, 0x2B,
	0x0B, 0x20, 0x26, 0x17, 0x59, 0x39, 0x20, 0x2E, 0x0D, 0x3A, 0x50, 0x3B,
	0x19, 0x29, 0x1F, 0x39, 0x06, 0x0A, 0x6D, 0x19, 0x1B, 0x3D, 0x3E, 0x69,
	0x5C, 0x38, 0x1E, 0x00, 0x2D, 0x39, 0x14, 0x57, 0x5E, 0x28, 0x0F, 0x58,
	0x28, 0x52, 0x7B, 0x5D, 0x53, 0x23, 0x53, 0x14, 0x2F, 0x18, 0x25, 0x04,
	0x23, 0x5C, 0x10, 0x2A, 0x00, 0x31, 0x2A, 0x4A, 0x08, 0x5D, 0x2E, 0x3C,
	0x2C, 0x5D, 0x1A, 0x76, 0x34, 0x09, 0x00, 0x18, 0x03, 0x16, 0x34, 0x03,
	0x08, 0x10, 0x1A, 0x00, 0x45, 0x2F, 0x37, 0x16, 0x0C, 0x5C, 0x58, 0x69,
	0x1B, 0x55, 0x0F, 0x21, 0x14, 0x1E, 0x0C, 0x19, 0x23, 0x7A, 0x04, 0x34,
	0x23, 0x0A, 0x0C, 0x09, 0x59, 0x07, 0x5F, 0x29, 0x15, 0x36, 0x56, 0x5E,
	0x15, 0x24, 0x19, 0x21, 0x5F, 0x06, 0x29, 0x2F, 0x00, 0x58, 0x11, 0x43,
	0x32, 0x1C, 0x1B, 0x2F, 0x3F, 0x23, 0x24, 0x06, 0x71, 0x39, 0x26, 0x2C,
	0x01, 0x72, 0x5E, 0x0E, 0x1B, 0x0F, 0x2F, 0x39, 0x06, 0x04, 0x33, 0x77,
	0x03, 0x17, 0x2C, 0x03, 0x17, 0x55, 0x27, 0x18, 0x22, 0x09, 0x1A, 0x02,
	0x3E, 0x22, 0x21, 0x0B, 0x0D, 0x0F, 0x23, 0x20, 0x3F, 0x17, 0x58, 0x5D,
	0x05, 0x19, 0x3B, 0x23, 0x3E, 0x1A, 0x05, 0x2D, 0x29, 0x5A, 0x72, 0x18,
	0x27, 0x5E, 0x58, 0x77, 0x0B, 0x35, 0x0F, 0x05, 0x03, 0x1E, 0x28, 0x1E,
	0x58, 0x1B, 0x5E, 0x4A, 0x3C, 0x1F, 0x0D, 0x19, 0x36, 0x0F, 0x01, 0x7B,
	0x28, 0x08, 0x5B, 0x3F, 0x32, 0x1B, 0x2B, 0x57, 0x29, 0x7B, 0x54, 0x2F,
	0x19, 0x44, 0x07, 0x5A, 0x15, 0x03, 0x3B, 0x16, 0x2E, 0x39, 0x18, 0x39,
	0x32, 0x39, 0x0E, 0x59, 0x24, 0x77, 0x00, 0x54, 0x2F, 0x31, 0x74, 0x38,
	0x51, 0x17, 0x12, 0x69, 0x58, 0x54, 0x2B, 0x32, 0x73, 0x3D, 0x1B, 0x03,
	0x04, 0x30, 0x39, 0x02, 0x2B, 0x59, 0x1B, 0x18, 0x20, 0x5D, 0x22, 0x0B,
	0x15, 0x26, 0x5F, 0x04, 0x04, 0x3D, 0x29, 0x41, 0x3C, 0x0A, 0x58, 0x30,
	0x5F, 0x3C, 0x2C, 0x2E, 0x06, 0x59, 0x2C, 0x72, 0x0B, 0x02, 0x18, 0x31,
	0x24, 0x2E, 0x35, 0x04, 0x0D, 0x73, 0x5C, 0x16, 0x5D, 0x27, 0x1A, 0x23,
	0x04, 0x17, 0x19, 0x77, 0x18, 0x57, 0x18, 0x2F, 0x13, 0x59, 0x52, 0x00,
	0x32, 0x29, 0x3C, 0x50, 0x06, 0x04, 0x21, 0x5A, 0x52, 0x3B, 0x3D, 0x06,
	0x1A, 0x34, 0x27, 0x09, 0x23, 0x1E, 0x17, 0x02, 0x44, 0x3B, 0x07, 0x38,
	0x1D, 0x3F, 0x6D, 0x29, 0x24, 0x00, 0x5E, 0x69, 0x3C, 0x35, 0x1D, 0x5D,
	0x2A, 0x00, 0x53, 0x0F, 0x06, 0x33, 0x2B, 0x13, 0x0C, 0x20, 0x0E, 0x01,
	0x06, 0x24, 0x1B, 0x0E, 0x43, 0x35, 0x1A, 0x0D, 0x2D, 0x5B, 0x56, 0x0C,
	0x13, 0x1A, 0x21, 0x18, 0x45, 0x5D, 0x38, 0x20, 0x27, 0x07, 0x28, 0x28,
	0x0F, 0x08, 0x07, 0x3F, 0x30, 0x43, 0x20, 0x36, 0x19, 0x69, 0x35, 0x54,
	0x58, 0x2D, 0x76, 0x5E, 0x25, 0x37, 0x2A, 0x24, 0x05, 0x19, 0x27, 0x08,
	0x10, 0x18, 0x10, 0x5B, 0x26, 0x70, 0x1A, 0x19, 0x28, 0x28, 0x0A, 0x38,
	0x00, 0x59, 0x44, 0x35, 0x5F, 0x22, 0x3B, 0x53, 0x00, 0x59, 0x0F, 0x2A,
	0x40, 0x12, 0x21, 0x20, 0x00, 0x39, 0x06, 0x5C, 0x0E, 0x5D, 0x0A, 0x25,
	0x38, 0x58, 0x04, 0x31, 0x20, 0x3B, 0x2D, 0x1E, 0x52, 0x3A, 0x3F, 0x50,
	0x18, 0x20, 0x04, 0x2D, 0x2C, 0x39, 0x5F, 0x30, 0x59, 0x58, 0x29, 0x3F,
	0x2A, 0x3F, 0x00, 0x08, 0x18, 0x16, 0x07, 0x2D, 0x39, 0x23, 0x0A, 0x5E,
	0x02, 0x3F, 0x2F, 0x38, 0x0E, 0x4A, 0x5D, 0x5D, 0x28, 0x58, 0x53, 0x08,
	0x3A, 0x36, 0x54, 0x15, 0x07, 0x5B, 0x38, 0x03, 0x4A, 0x0F, 0x1E, 0x27,
	0x25, 0x09, 0x21, 0x2C, 0x05, 0x39, 0x58, 0x2A, 0x12, 0x7A, 0x5B, 0x1B,
	0x2F, 0x03, 0x74, 0x21, 0x09, 0x58, 0x23, 0x73, 0x27, 0x32, 0x03, 0x05,
	0x0D, 0x36, 0x38, 0x0D, 0x13, 0x2D, 0x0A, 0x06, 0x18, 0x04, 0x1A, 0x18,
	0x57, 0x24, 0x2D, 0x2C, 0x36, 0x28, 0x41, 0x00, 0x16, 0x38, 0x15, 0x3E,
	0x18, 0x37, 0x1B, 0x11, 0x58, 0x03, 0x12, 0x26, 0x17, 0x06, 0x21, 0x10,
	0x1A, 0x4A, 0x3F, 0x0C, 0x03, 0x5C, 0x14, 0x2A, 0x0E, 0x31, 0x54, 0x4A,
	0x39, 0x0C, 0x2F, 0x5F, 0x0C, 0x0C, 0x00, 0x2C, 0x04, 0x4A, 0x41, 0x3A,
	0x0F, 0x5E, 0x50, 0x00, 0x20, 0x3A, 0x0E, 0x25, 0x09, 0x2C, 0x26, 0x47,
	0x59, 0x2F, 0x5F, 0x7B, 0x5E, 0x57, 0x04, 0x01, 0x12, 0x55, 0x0B, 0x45,
	0x2F, 0x7B, 0x1F, 0x08, 0x2F, 0x59, 0x01, 0x0B, 0x2E, 0x3A, 0x1D, 0x23,
	0x5B, 0x02, 0x08, 0x2E, 0x74, 0x36, 0x0A, 0x3B, 0x5D, 0x36, 0x35, 0x30,
	0x01, 0x58, 0x0E, 0x26, 0x32, 0x29, 0x03, 0x7A, 0x2A, 0x17, 0x0F, 0x29,
	0x26, 0x07, 0x0E, 0x2D, 0x11, 0x35, 0x54, 0x52, 0x3B, 0x2E, 0x3B, 0x09,
	0x16, 0x1E, 0x53, 0x20, 0x38, 0x36, 0x17, 0x5D, 0x00, 0x04, 0x2C, 0x00,
	0x21, 0x1B, 0x03, 0x14, 0x5D, 0x0C, 0x01, 0x1C, 0x38, 0x26, 0x1B, 0x0F,
	0x21, 0x0D, 0x1D, 0x19, 0x7A, 0x1A, 0x15, 0x17, 0x5D, 0x28, 0x3A, 0x4E,
	0x01, 0x21, 0x13, 0x1B, 0x05, 0x0A, 0x5A, 0x0D, 0x09, 0x16, 0x0D, 0x27,
	0x72, 0x2B, 0x1B, 0x2A, 0x5B, 0x0F, 0x0B, 0x0C, 0x5D, 0x29, 0x01, 0x3D,
	0x35, 0x3B, 0x58, 0x0B, 0x25, 0x18, 0x1C, 0x27, 0x70, 0x29, 0x56, 0x1B,
	0x28, 0x0A, 0x38, 0x27, 0x3A, 0x40, 0x77, 0x26, 0x23, 0x37, 0x08, 0x2C,
	0x0D, 0x3B, 0x59, 0x58, 0x14, 0x35, 0x06, 0x1E, 0x07, 0x2C, 0x1E, 0x23,
	0x57, 0x39, 0x71, 0x3E, 0x58, 0x36, 0x2D, 0x3A, 0x3B, 0x2E, 0x1C, 0x07,
	0x2F, 0x5E, 0x20, 0x24, 0x1E, 0x72, 0x1E, 0x18, 0x19, 0x22, 0x31, 0x5F,
	0x38, 0x0F, 0x2C, 0x13, 0x03, 0x57, 0x1D, 0x04, 0x18, 0x59, 0x57, 0x57,
	0x20, 0x10, 0x03, 0x2D, 0x5F, 0x12, 0x77, 0x09, 0x22, 0x5F, 0x2F, 0x70,
	0x5C, 0x33, 0x3B, 0x32, 0x05, 0x01, 0x03, 0x57, 0x2E, 0x11, 0x0E, 0x2A,
	0x1F, 0x08, 0x6D, 0x19, 0x33, 0x03, 0x3D, 0x73, 0x22, 0x35, 0x36, 0x44,
	0x0D, 0x38, 0x31, 0x0F, 0x13, 0x7B, 0x28, 0x16, 0x56, 0x1A, 0x38, 0x5C,
	0x18, 0x22, 0x1C, 0x03, 0x36, 0x06, 0x20, 0x2A, 0x26, 0x07, 0x54, 0x3F,
	0x40, 0x03, 0x19, 0x52, 0x01, 0x32, 0x09, 0x0D, 0x0C, 0x0C, 0x5F, 0x26,
	0x24, 0x16, 0x21, 0x5C, 0x13, 0x3D, 0x03, 0x39, 0x12, 0x25, 0x21, 0x51,
	0x22, 0x3A, 0x06, 0x08, 0x18, 0x39, 0x1E, 0x7A, 0x29, 0x06, 0x57, 0x3D,
	0x26, 0x28, 0x59, 0x25, 0x1A, 0x08, 0x1F, 0x33, 0x57, 0x05, 0x26, 0x27,
	0x52, 0x1D, 0x23, 0x26, 0x3E, 0x31, 0x56, 0x1E, 0x12, 0x1A, 0x09, 0x0F,
	0x0E, 0x0C, 0x55, 0x55, 0x34, 0x2A, 0x31, 0x0E, 0x4A, 0x2A, 0x26, 0x20,
	0x15, 0x3B, 0x3D, 0x53, 0x34, 0x1B, 0x07, 0x27, 0x53, 0x04, 0x07, 0x0B,
	0x05, 0x09, 0x11, 0x19, 0x19, 0x2A, 0x2A, 0x3B, 0x2E, 0x2A, 0x28, 0x53,
	0x13, 0x26, 0x2B, 0x5D, 0x1A, 0x20, 0x0D, 0x30, 0x04, 0x0C, 0x37, 0x47,
	0x12, 0x2F, 0x20, 0x12, 0x5E, 0x10, 0x07, 0x44, 0x75, 0x21, 0x2B, 0x3C,
	0x40, 0x2D, 0x05, 0x18, 0x3B, 0x5E, 0x07, 0x58, 0x1B, 0x17, 0x24, 0x73,
	0x04, 0x4E, 0x56, 0x32, 0x10, 0x47, 0x33, 0x57, 0x12, 0x01, 0x1B, 0x23,
	0x0F, 0x44, 0x1A, 0x1A, 0x2C, 0x1F, 0x02, 0x0E, 0x08, 0x51, 0x38, 0x06,
	0x76, 0x5B, 0x0C, 0x23, 0x03, 0x18, 0x0B, 0x59, 0x23, 0x1C, 0x16, 0x55,
	0x29, 0x59, 0x40, 0x11, 0x43, 0x57, 0x23, 0x2C, 0x20, 0x27, 0x0D, 0x14,
	0x3A, 0x75, 0x24, 0x19, 0x08, 0x5C, 0x28, 0x0A, 0x16, 0x57, 0x2A, 0x71,
	0x08, 0x1B, 0x03, 0x2D, 0x69, 0x2A, 0x0B, 0x56, 0x2A, 0x12, 0x1F, 0x10,
	0x0F, 0x3B, 0x33, 0x01, 0x0C, 0x3D, 0x1C, 0x31, 0x2F, 0x25, 0x08, 0x59,
	0x16, 0x5E, 0x1B, 0x26, 0x5B, 0x0F, 0x08, 0x24, 0x5E, 0x3D, 0x37, 0x0B,
	0x22, 0x5A, 0x00, 0x06, 0x15, 0x08, 0x28, 0x58, 0x35, 0x5F, 0x2C, 0x3B,
	0x0F, 0x0D, 0x38, 0x0E, 0x07, 0x53, 0x31, 0x14, 0x57, 0x19, 0x19, 0x07,
	0x58, 0x0E, 0x16, 0x5D, 0x21, 0x3E, 0x06, 0x41, 0x1E, 0x03, 0x2B, 0x0F,
	0x23, 0x5B, 0x28, 0x24, 0x59, 0x26, 0x3D, 0x0B, 0x25, 0x50, 0x24, 0x1C,
	0x08, 0x3D, 0x27, 0x36, 0x01, 0x38, 0x16, 0x05, 0x5C, 0x2D, 0x2A, 0x3C,
	0x55, 0x07, 0x2A, 0x12, 0x05, 0x0E, 0x26, 0x2A, 0x7B, 0x0B, 0x18, 0x05,
	0x0C, 0x2D, 0x43, 0x39, 0x2F, 0x5A, 0x08, 0x0F, 0x54, 0x1F, 0x24, 0x36,
	0x02, 0x29, 0x1F, 0x59, 0x2E, 0x0A, 0x2F, 0x1F, 0x2A, 0x70, 0x5F, 0x0D,
	0x0B, 0x29, 0x2D, 0x05, 0x36, 0x14, 0x00, 0x34, 0x43, 0x19, 0x17, 0x11,
	0x2E, 0x38, 0x2C, 0x1B, 0x28, 0x20, 0x08, 0x18, 0x1E, 0x1D, 0x38, 0x0F,
	0x02, 0x3D, 0x18, 0x0A, 0x55, 0x52, 0x2D, 0x53, 0x1A, 0x54, 0x2C, 0x18,
	0x3B, 0x21, 0x0D, 0x19, 0x5F, 0x2F, 0x12, 0x24, 0x16, 0x21, 0x59, 0x2B,
	0x1C, 0x00, 0x36, 0x5F, 0x26, 0x1D, 0x09, 0x57, 0x3B, 0x2B, 0x2A, 0x03,
	0x1E, 0x3F, 0x03, 0x20, 0x58, 0x59, 0x26, 0x0B, 0x1A, 0x34, 0x45, 0x28,
	0x17, 0x38, 0x55, 0x0C, 0x02, 0x33, 0x01, 0x39, 0x3B, 0x3D, 0x3B, 0x2D,
	0x57, 0x38, 0x2C, 0x31, 0x58, 0x0F, 0x38, 0x0D, 0x00, 0x1A, 0x0A, 0x06,
	0x39, 0x0F, 0x1F, 0x55, 0x08, 0x25, 0x35, 0x3C, 0x08, 0x16, 0x33, 0x27,
	0x04, 0x59, 0x1E, 0x07, 0x38, 0x01, 0x50, 0x3E, 0x5D, 0x0D, 0x00, 0x31,
	0x19, 0x24, 0x1B, 0x39, 0x2C, 0x5B, 0x1A, 0x35, 0x06, 0x18, 0x45, 0x0C,
	0x2A, 0x36, 0x04, 0x58, 0x22, 0x1B, 0x5E, 0x37, 0x07, 0x08, 0x08, 0x5D,
	0x08, 0x20, 0x3A, 0x37, 0x09, 0x20, 0x18, 0x24, 0x28, 0x47, 0x28, 0x08,
	0x09, 0x23, 0x26, 0x07, 0x05, 0x1C, 0x29, 0x08, 0x50, 0x06, 0x1C, 0x05,
	0x43, 0x11, 0x1C, 0x1F, 0x01, 0x5F, 0x56, 0x22, 0x44, 0x0E, 0x5A, 0x0C,
	0x06, 0x52, 0x26, 0x1E, 0x58, 0x3B, 0x31, 0x25, 0x1A, 0x35, 0x18, 0x03,
	0x28, 0x3B, 0x53, 0x5D, 0x0A, 0x0A, 0x15, 0x05, 0x1C, 0x52, 0x2F, 0x1D,
	0x54, 0x19, 0x04, 0x17, 0x1A, 0x0B, 0x1D, 0x25, 0x72, 0x24, 0x06, 0x24,
	0x05, 0x2E, 0x02, 0x16, 0x18, 0x1B, 0x2D, 0x3D, 0x51, 0x1E, 0x2E, 0x14,
	0x5E, 0x27, 0x5F, 0x52, 0x05, 0x36, 0x0E, 0x22, 0x0D, 0x0C, 0x5F, 0x36,
	0x0C, 0x05, 0x69, 0x15, 0x0F, 0x0C, 0x59, 0x21, 0x34, 0x11, 0x04, 0x0F,
	0x75, 0x21, 0x10, 0x59, 0x32, 0x3B, 0x19, 0x3B, 0x41, 0x1E, 0x34, 0x00,
	0x13, 0x37, 0x27, 0x75, 0x2D, 0x0C, 0x3F, 0x07, 0x71, 0x03, 0x27, 0x41,
	0x21, 0x09, 0x26, 0x05, 0x38, 0x1B, 0x03, 0x2B, 0x00, 0x5B, 0x11, 0x77,
	0x5C, 0x27, 0x34, 0x18, 0x27, 0x00, 0x2A, 0x07, 0x5E, 0x04, 0x5E, 0x34,
	0x07, 0x2C, 0x1B, 0x39, 0x13, 0x1A, 0x5E, 0x2C, 0x3E, 0x23, 0x1C, 0x33,
	0x2E, 0x22, 0x0E, 0x57, 0x22, 0x21, 0x2A, 0x05, 0x17, 0x01, 0x10, 0x35,
	0x33, 0x41, 0x0F, 0x13, 0x24, 0x32, 0x22, 0x0A, 0x00, 0x1F, 0x18, 0x3A,
	0x3C, 0x76, 0x2B, 0x05, 0x59, 0x25, 0x7A, 0x0D, 0x54, 0x04, 0x00, 0x10,
	0x54, 0x52, 0x34, 0x25, 0x28, 0x24, 0x0F, 0x1C, 0x5C, 0x00, 0x1A, 0x12,
	0x41, 0x44, 0x26, 0x5E, 0x03, 0x39, 0x18, 0x75, 0x3C, 0x56, 0x0B, 0x38,
	0x09, 0x21, 0x0E, 0x57, 0x0C, 0x23, 0x04, 0x23, 0x2A, 0x3F, 0x27, 0x55,
	0x34, 0x3F, 0x1D, 0x38, 0x2A, 0x54, 0x0F, 0x21, 0x6D, 0x39, 0x35, 0x36,
	0x2A, 0x18, 0x5F, 0x2F, 0x3B, 0x1E, 0x0F, 0x35, 0x00, 0x34, 0x26, 0x71,
	0x58, 0x52, 0x09, 0x53, 0x29, 0x5E, 0x09, 0x00, 0x1D, 0x3B, 0x20, 0x33,
	0x34, 0x1D, 0x2E, 0x38, 0x59, 0x20, 0x12, 0x01, 0x3A, 0x20, 0x3F, 0x26,
	0x0A, 0x47, 0x2E, 0x24, 0x32, 0x04, 0x27, 0x32, 0x1E, 0x3D, 0x0A, 0x1B,
	0x39, 0x27, 0x29, 0x2C, 0x05, 0x31, 0x22, 0x1E, 0x71, 0x1B, 0x2D, 0x3A,
	0x0F, 0x2D, 0x15, 0x06, 0x2C, 0x3A, 0x38, 0x5E, 0x25, 0x56, 0x25, 0x73,
	0x28, 0x23, 0x2A, 0x3B, 0x11, 0x08, 0x39, 0x19, 0x2F, 0x25, 0x0E, 0x4A,
	0x36, 0x03, 0x12, 0x03, 0x35, 0x16, 0x1D, 0x2B, 0x1F, 0x03, 0x19, 0x2F,
	0x28, 0x0D, 0x25, 0x17, 0x00, 0x0D, 0x02, 0x04, 0x14, 0x0A, 0x01, 0x2F,
	0x18, 0x16, 0x3C, 0x00, 0x5A, 0x0B, 0x0F, 0x00, 0x32, 0x2E, 0x12, 0x5D,
	0x00, 0x71, 0x2F, 0x20, 0x0A, 0x0A, 0x2B, 0x5B, 0x23, 0x2B, 0x0A, 0x14,
	0x5C, 0x32, 0x3D, 0x33, 0x33, 0x0E, 0x52, 0x2F, 0x0F, 0x03, 0x04, 0x4A,
	0x5E, 0x2D, 0x76, 0x47, 0x19, 0x23, 0x26, 0x6D, 0x3A, 0x52, 0x3F, 0x52,
	0x29, 0x1B, 0x54, 0x25, 0x1C, 0x3B, 0x47, 0x22, 0x5C, 0x5D, 0x32, 0x24,
	0x2F, 0x26, 0x04, 0x2F, 0x2A, 0x56, 0x04, 0x53, 0x04, 0x0A, 0x09, 0x3A,
	0x0E, 0x21, 0x35, 0x2C, 0x0B, 0x03, 0x3A, 0x21, 0x22, 0x0A, 0x0C, 0x2F,
	0x43, 0x18, 0x3E, 0x3B, 0x74, 0x3F, 0x33, 0x02, 0x5F, 0x0D, 0x3D, 0x15,
	0x5B, 0x23, 0x3B, 0x0D, 0x20, 0x01, 0x52, 0x09, 0x43, 0x14, 0x23, 0x1F,
	0x16, 0x21, 0x1B, 0x0F, 0x5E, 0x06, 0x36, 0x34, 0x21, 0x26, 0x11, 0x3F,
	0x24, 0x29, 0x07, 0x29, 0x16, 0x14, 0x14, 0x06, 0x1B, 0x29, 0x0E, 0x3B,
	0x1D, 0x71, 0x3E, 0x0F, 0x3D, 0x26, 0x7A, 0x58, 0x28, 0x1D, 0x13, 0x33,
	0x25, 0x2F, 0x1F, 0x20, 0x73, 0x16, 0x2E, 0x25, 0x0D, 0x75, 0x21, 0x13,
	0x06, 0x0E, 0x2F, 0x58, 0x12, 0x0C, 0x1C, 0x04, 0x23, 0x27, 0x2B, 0x12,
	0x03, 0x27, 0x02, 0x27, 0x2F, 0x03, 0x2E, 0x4A, 0x3B, 0x12, 0x75, 0x14,
	0x0E, 0x1B, 0x2D, 0x20, 0x5C, 0x2A, 0x5C, 0x3D, 0x7B, 0x1B, 0x14, 0x1E,
	0x33, 0x18, 0x58, 0x0F, 0x2B, 0x5B, 0x2B, 0x5D, 0x32, 0x17, 0x32, 0x23,
	0x38, 0x06, 0x0A, 0x3C, 0x0B, 0x21, 0x0F, 0x5B, 0x02, 0x15, 0x29, 0x58,
	0x19, 0x40, 0x18, 0x1D, 0x51, 0x19, 0x1D, 0x37, 0x09, 0x4E, 0x3A, 0x5B,
	0x01, 0x47, 0x19, 0x3C, 0x25, 0x69, 0x01, 0x23, 0x24, 0x0A, 0x16, 0x5F,
	0x14, 0x25, 0x2A, 0x34, 0x05, 0x50, 0x57, 0x1C, 0x71, 0x39, 0x3B, 0x1E,
	0x27, 0x71, 0x2A, 0x0A, 0x45, 0x24, 0x23, 0x54, 0x34, 0x27, 0x3D, 0x23,
	0x08, 0x50, 0x5B, 0x13, 0x04, 0x5B, 0x03, 0x41, 0x59, 0x3A, 0x09, 0x20,
	0x5D, 0x23, 0x2A, 0x2B, 0x05, 0x3E, 0x00, 0x0F, 0x59, 0x22, 0x21, 0x1C,
	0x09, 0x08, 0x2E, 0x16, 0x22, 0x37, 0x04, 0x50, 0x09, 0x2D, 0x7A, 0x1F,
	0x30, 0x3E, 0x26, 0x35, 0x1B, 0x08, 0x45, 0x44, 0x37, 0x3A, 0x28, 0x00,
	0x1E, 0x12, 0x0F, 0x35, 0x16, 0x1D, 0x11, 0x5C, 0x36, 0x3A, 0x31, 0x12,
	0x23, 0x02, 0x1A, 0x06, 0x70, 0x38, 0x32, 0x5B, 0x21, 0x77, 0x2F, 0x33,
	0x36, 0x3C, 0x77, 0x39, 0x53, 0x45, 0x1B, 0x73, 0x14, 0x2A, 0x21, 0x3E,
	0x74, 0x14, 0x2C, 0x59, 0x5E, 0x0D, 0x5E, 0x2E, 0x5B, 0x28, 0x14, 0x5F,
	0x18, 0x25, 0x1E, 0x0B, 0x59, 0x2A, 0x38, 0x5B, 0x3B, 0x3C, 0x12, 0x1D,
	0x00, 0x2F, 0x0A, 0x14, 0x05, 0x2F, 0x21, 0x1A, 0x0A, 0x1E, 0x0D, 0x27,
	0x25, 0x00, 0x56, 0x04, 0x29, 0x1C, 0x07, 0x38, 0x22, 0x27, 0x47, 0x36,
	0x3D, 0x2D, 0x76, 0x19, 0x54, 0x18, 0x33, 0x06, 0x3C, 0x2B, 0x21, 0x3C,
	0x26, 0x14, 0x39, 0x22, 0x28, 0x7B, 0x23, 0x27, 0x1F, 0x12, 0x08, 0x0A,
	0x58, 0x2C, 0x53, 0x00, 0x05, 0x2E, 0x01, 0x39, 0x33, 0x39, 0x17, 0x39,
	0x22, 0x12, 0x3E, 0x24, 0x5F, 0x59, 0x0C, 0x1C, 0x57, 0x0F, 0x29, 0x73,
	0x0E, 0x55, 0x5D, 0x5D, 0x23, 0x5C, 0x34, 0x5B, 0x52, 0x20, 0x5A, 0x07,
	0x57, 0x39, 0x07, 0x47, 0x27, 0x2B, 0x2D, 0x17, 0x3B, 0x20, 0x5C, 0x0F,
	0x2D, 0x59, 0x4E, 0x05, 0x33, 0x17, 0x29, 0x13, 0x05, 0x3A, 0x04, 0x2B,
	0x1B, 0x0B, 0x0A, 0x2B, 0x19, 0x0A, 0x2A, 0x2F, 0x2F, 0x3D, 0x06, 0x08,
	0x02, 0x14, 0x19, 0x0B, 0x5A, 0x1E, 0x1A, 0x3E, 0x58, 0x3A, 0x07, 0x13,
	0x3D, 0x04, 0x1A, 0x3F, 0x18, 0x43, 0x08, 0x22, 0x52, 0x1A, 0x2A, 0x10,
	0x58, 0x52, 0x12, 0x1F, 0x26, 0x2D, 0x1D, 0x09, 0x3E, 0x59, 0x22, 0x5F,
	0x2E, 0x18, 0x58, 0x0D, 0x04, 0x1A, 0x22, 0x02, 0x24, 0x38, 0x32, 0x2F,
	0x09, 0x14, 0x05, 0x6D, 0x36, 0x57, 0x1D, 0x59, 0x77, 0x14, 0x15, 0x01,
	0x09, 0x21, 0x5B, 0x26, 0x18, 0x2D, 0x77, 0x0D, 0x52, 0x1C, 0x3D, 0x20,
	0x18, 0x35, 0x00, 0x2F, 0x00, 0x2F, 0x10, 0x3A, 0x13, 0x18, 0x1E, 0x25,
	0x14, 0x06, 0x14, 0x14, 0x34, 0x5D, 0x3C, 0x15, 0x07, 0x11, 0x04, 0x28,
	0x6D, 0x24, 0x38, 0x5A, 0x31, 0x11, 0x2F, 0x09, 0x28, 0x03, 0x75, 0x16,
	0x27, 0x39, 0x11, 0x0F, 0x59, 0x4E, 0x41, 0x01, 0x2F, 0x2D, 0x36, 0x5D,
	0x3F, 0x07, 0x2D, 0x56, 0x3F, 0x1E, 0x0F, 0x18, 0x57, 0x03, 0x12, 0x7A,
	0x43, 0x58, 0x1D, 0x38, 0x0C, 0x55, 0x57, 0x5A, 0x1D, 0x0C, 0x0F, 0x08,
	0x0B, 0x39, 0x73, 0x14, 0x57, 0x34, 0x07, 0x0B, 0x34, 0x0A, 0x1F, 0x23,
	0x27, 0x08, 0x57, 0x14, 0x21, 0x15, 0x0D, 0x04, 0x34, 0x1F, 0x04, 0x43,
	0x36, 0x2D, 0x52, 0x76, 0x02, 0x14, 0x03, 0x5F, 0x30, 0x06, 0x04, 0x04,
	0x52, 0x0E, 0x54, 0x38, 0x57, 0x5A, 0x14, 0x22, 0x32, 0x5C, 0x1A, 0x08,
	0x19, 0x18, 0x45, 0x40, 0x11, 0x21, 0x4E, 0x56, 0x5F, 0x0D, 0x1E, 0x52,
	0x25, 0x1B, 0x33, 0x3C, 0x59, 0x2D, 0x18, 0x35, 0x2F, 0x30, 0x3C, 0x3E,
	0x23, 0x08, 0x06, 0x41, 0x5C, 0x27, 0x34, 0x2D, 0x0F, 0x18, 0x2B, 0x1A,
	0x07, 0x29, 0x08, 0x36, 0x47, 0x3B, 0x20, 0x3A, 0x75, 0x47, 0x19, 0x3B,
	0x59, 0x13, 0x1A, 0x29, 0x20, 0x1C, 0x08, 0x5F, 0x27, 0x03, 0x1D, 0x6D,
	0x23, 0x13, 0x5A, 0x13, 0x2D, 0x19, 0x4A, 0x5F, 0x5F, 0x75, 0x55, 0x35,
	0x5E, 0x5A, 0x05, 0x02, 0x24, 0x01, 0x23, 0x7B, 0x55, 0x10, 0x21, 0x39,
	0x1A, 0x36, 0x4A, 0x23, 0x18, 0x17, 0x3A, 0x2C, 0x14, 0x5D, 0x34, 0x2B,
	0x24, 0x38, 0x01, 0x7A, 0x3E, 0x02, 0x23, 0x1C, 0x24, 0x01, 0x2C, 0x01,
	0x08, 0x18, 0x2D, 0x1B, 0x20, 0x08, 0x2A, 0x2E, 0x35, 0x02, 0x3D, 0x16,
	0x23, 0x31, 0x2A, 0x3D, 0x2D, 0x1A, 0x16, 0x1B, 0x08, 0x1B, 0x47, 0x32,
	0x19, 0x5B, 0x71, 0x02, 0x28, 0x41, 0x39, 0x2C, 0x2D, 0x25, 0x08, 0x3B,
	0x69, 0x0D, 0x16, 0x03, 0x32, 0x32, 0x2B, 0x34, 0x5A, 0x44, 0x75, 0x1E,
	0x2B, 0x02, 0x2E, 0x69, 0x38, 0x59, 0x1A, 0x5D, 0x0F, 0x3F, 0x38, 0x22,
	0x0C, 0x0E, 0x2E, 0x0E, 0x2B, 0x2E, 0x28, 0x26, 0x56, 0x5D, 0x44, 0x0A,
	0x5B, 0x00, 0x2B, 0x22, 0x24, 0x1B, 0x14, 0x0D, 0x02, 0x32, 0x08, 0x16,
	0x0D, 0x0E, 0x21, 0x34, 0x16, 0x2F, 0x1C, 0x05, 0x55, 0x14, 0x00, 0x0D,
	0x18, 0x5C, 0x22, 0x1C, 0x5F, 0x1B, 0x3C, 0x57, 0x3B, 0x2E, 0x2B, 0x20,
	0x56, 0x07, 0x03, 0x1A, 0x09, 0x26, 0x05, 0x2F, 0x06, 0x1F, 0x0D, 0x16,
	0x27, 0x36, 0x0B, 0x29, 0x29, 0x52, 0x01, 0x5B, 0x2D, 0x38, 0x0D, 0x72,
	0x15, 0x27, 0x2B, 0x05, 0x7A, 0x59, 0x16, 0x19, 0x1D, 0x35, 0x14, 0x55,
	0x26, 0x39, 0x73, 0x01, 0x23, 0x39, 0x28, 0x70, 0x3A, 0x04, 0x20, 0x29,
	0x74, 0x47, 0x13, 0x24, 0x1E, 0x08, 0x18, 0x58, 0x39, 0x32, 0x73, 0x09,
	0x51, 0x16, 0x02, 0x20, 0x24, 0x30, 0x45, 0x01, 0x36, 0x26, 0x2C, 0x3B,
	0x5F, 0x35, 0x39, 0x55, 0x23, 0x3F, 0x06, 0x3E, 0x3B, 0x03, 0x28, 0x74,
	0x5D, 0x52, 0x2F, 0x21, 0x17, 0x23, 0x29, 0x58, 0x0A, 0x34, 0x20, 0x13,
	0x00, 0x5D, 0x1B, 0x24, 0x17, 0x58, 0x0A, 0x23, 0x5A, 0x35, 0x39, 0x44,
	0x07, 0x05, 0x0A, 0x26, 0x2A, 0x14, 0x05, 0x11, 0x25, 0x5D, 0x34, 0x0E,
	0x57, 0x0F, 0x27, 0x23, 0x0A, 0x0F, 0x27, 0x19, 0x38, 0x3C, 0x23, 0x0F,
	0x05, 0x0D, 0x24, 0x00, 0x41, 0x0A, 0x2A, 0x58, 0x11, 0x23, 0x5D, 0x01,
	0x0F, 0x12, 0x26, 0x5A, 0x77, 0x2E, 0x0B, 0x0F, 0x2C, 0x05, 0x5F, 0x4A,
	0x23, 0x0F, 0x20, 0x54, 0x2E, 0x58, 0x11, 0x77, 0x05, 0x37, 0x04, 0x06,
	0x07, 0x5A, 0x38, 0x18, 0x53, 0x0C, 0x55, 0x2C, 0x16, 0x19, 0x0F, 0x21,
	0x31, 0x20, 0x0A, 0x16, 0x1A, 0x2E, 0x3E, 0x39, 0x09, 0x5C, 0x33, 0x26,
	0x26, 0x13, 0x0E, 0x59, 0x27, 0x3C, 0x1A, 0x1F, 0x15, 0x00, 0x1D, 0x70,
	0x3F, 0x0A, 0x22, 0x03, 0x20, 0x1E, 0x15, 0x02, 0x0F, 0x26, 0x2A, 0x20,
	0x14, 0x5A, 0x30, 0x24, 0x4E, 0x58, 0x28, 0x34, 0x2A, 0x16, 0x0F, 0x02,
	0x36, 0x34, 0x0E, 0x5E, 0x1E, 0x73, 0x36, 0x58, 0x2D, 0x2F, 0x32, 0x39,
	0x0B, 0x22, 0x0F, 0x31, 0x2E, 0x06, 0x36, 0x01, 0x3B, 0x1C, 0x22, 0x03,
	0x1B, 0x7B, 0x1E, 0x0D, 0x20, 0x0E, 0x09, 0x26, 0x04, 0x00, 0x1D, 0x05,
	0x3C, 0x15, 0x1B, 0x2A, 0x0C, 0x0D, 0x20, 0x07, 0x33, 0x70, 0x34, 0x52,
	0x26, 0x23, 0x0B, 0x07, 0x0B, 0x08, 0x22, 0x2F, 0x28, 0x3B, 0x22, 0x00,
	0x03, 0x47, 0x0E, 0x5B, 0x13, 0x75, 0x24, 0x22, 0x3F, 0x20, 0x38, 0x3D,
	0x33, 0x37, 0x1E, 0x0E, 0x03, 0x04, 0x2B, 0x44, 0x01, 0x29, 0x53, 0x1F,
	0x44, 0x26, 0x06, 0x16, 0x17, 0x11, 0x05, 0x5F, 0x26, 0x16, 0x59, 0x07,
	0x23, 0x2C, 0x1F, 0x5B, 0x76, 0x0E, 0x57, 0x37, 0x0E, 0x3A, 0x03, 0x12,
	0x02, 0x02, 0x00, 0x5E, 0x39, 0x5A, 0x1B, 0x34, 0x59, 0x4A, 0x5E, 0x2D,
	0x74, 0x0E, 0x11, 0x39, 0x44, 0x23, 0x3D, 0x53, 0x28, 0x2C, 0x09, 0x02,
	0x56, 0x00, 0x53, 0x77, 0x1E, 0x14, 0x20, 0x20, 0x0D, 0x47, 0x18, 0x00,
	0x1B, 0x2D, 0x23, 0x2E, 0x1E, 0x40, 0x2A, 0x27, 0x02, 0x00, 0x06, 0x0D,
	0x54, 0x55, 0x26, 0x52, 0x14, 0x1D, 0x50, 0x28, 0x33, 0x36, 0x27, 0x59,
	0x36, 0x3D, 0x12, 0x22, 0x2E, 0x1B, 0x0F, 0x00, 0x3F, 0x33, 0x26, 0x3F,
	0x10, 0x3B, 0x4E, 0x1F, 0x1A, 0x29, 0x5D, 0x28, 0x41, 0x5D, 0x18, 0x3C,
	0x0F, 0x2F, 0x2A, 0x08, 0x18, 0x17, 0x26, 0x0A, 0x1B, 0x36, 0x07, 0x0A,
	0x2E, 0x2D, 0x5F, 0x17, 0x28, 0x3F, 0x24, 0x43, 0x30, 0x5D, 0x1C, 0x34,
	0x0D, 0x18, 0x21, 0x26, 0x6D, 0x5A, 0x57, 0x1C, 0x1A, 0x38, 0x07, 0x57,
	0x17, 0x05, 0x73, 0x0E, 0x2C, 0x39, 0x02, 0x2F, 0x1E, 0x11, 0x0F, 0x3A,
	0x2D, 0x16, 0x02, 0x0C, 0x02, 0x00, 0x04, 0x10, 0x04, 0x24, 0x00, 0x06,
	0x05, 0x03, 0x58, 0x25, 0x20, 0x0D, 0x27, 0x1E, 0x36, 0x19, 0x09, 0x2F,
	0x24, 0x29, 0x18, 0x51, 0x3C, 0x0C, 0x38, 0x35, 0x51, 0x27, 0x06, 0x26,
	0x5C, 0x0E, 0x2C, 0x25, 0x30, 0x1F, 0x03, 0x38, 0x00, 0x36, 0x0A, 0x38,
	0x29, 0x1C, 0x18, 0x34, 0x55, 0x23, 0x58, 0x12, 0x1C, 0x51, 0x21, 0x3C,
	0x37, 0x05, 0x0E, 0x25, 0x39, 0x20, 0x54, 0x07, 0x39, 0x01, 0x71, 0x01,
	0x55, 0x25, 0x2C, 0x70, 0x2A, 0x15, 0x00, 0x03, 0x14, 0x59, 0x2C, 0x0D,
	0x29, 0x16, 0x3D, 0x4E, 0x45, 0x0A, 0x25, 0x08, 0x0D, 0x0B, 0x5D, 0x1B,
	0x20, 0x33, 0x5B, 0x09, 0x71, 0x3E, 0x56, 0x0F, 0x5E, 0x27, 0x2B, 0x07,
	0x59, 0x18, 0x7B, 0x14, 0x35, 0x38, 0x20, 0x71, 0x43, 0x10, 0x06, 0x44,
	0x0E, 0x58, 0x29, 0x0F, 0x3C, 0x07, 0x1A, 0x24, 0x56, 0x5A, 0x29, 0x00,
	0x27, 0x39, 0x3A, 0x25, 0x3B, 0x12, 0x1F, 0x20, 0x24, 0x2F, 0x15, 0x3C,
	0x3C, 0x35, 0x5E, 0x12, 0x24, 0x38, 0x1A, 0x00, 0x13, 0x09, 0x1A, 0x09,
	0x3F, 0x02, 0x1E, 0x24, 0x35, 0x59, 0x06, 0x05, 0x1F, 0x15, 0x0B, 0x17,
	0x03, 0x3A, 0x0F, 0x3F, 0x17, 0x25, 0x06, 0x06, 0x0D, 0x0B, 0x2A, 0x44,
	0x25, 0x38, 0x37, 0x09, 0x2F, 0x2A, 0x38, 0x27, 0x5C, 0x52, 0x16, 0x2D,
	0x36, 0x2C, 0x5C, 0x27, 0x2B, 0x23, 0x08, 0x3B, 0x7A, 0x47, 0x4E, 0x04,
	0x1B, 0x7B, 0x3B, 0x2F, 0x41, 0x44, 0x24, 0x58, 0x57, 0x0C, 0x5B, 0x20,
	0x5E, 0x12, 0x38, 0x3B, 0x2E, 0x5E, 0x4E, 0x3F, 0x44, 0x73, 0x5F, 0x59,
	0x20, 0x2C, 0x09, 0x20, 0x54, 0x2A, 0x3D, 0x7B, 0x18, 0x51, 0x2B, 0x27,
	0x36, 0x54, 0x23, 0x1A, 0x59, 0x11, 0x1E, 0x22, 0x2F, 0x21, 0x34, 0x05,
	0x2D, 0x01, 0x18, 0x0C, 0x07, 0x2C, 0x21, 0x5F, 0x2D, 0x5E, 0x12, 0x5D,
	0x0F, 0x2D, 0x05, 0x1B, 0x03, 0x29, 0x0D, 0x5F, 0x4E, 0x06, 0x3F, 0x34,
	0x3D, 0x2C, 0x21, 0x26, 0x10, 0x21, 0x0C, 0x28, 0x3B, 0x1B, 0x29, 0x38,
	0x5B, 0x5D, 0x15, 0x35, 0x51, 0x04, 0x32, 0x13, 0x2E, 0x52, 0x2F, 0x0D,
	0x76, 0x06, 0x35, 0x28, 0x40, 0x00, 0x39, 0x2E, 0x07, 0x3A, 0x21, 0x21,
	0x2B, 0x03, 0x26, 0x03, 0x14, 0x59, 0x2D, 0x02, 0x24, 0x01, 0x2D, 0x09,
	0x38, 0x1A, 0x29, 0x38, 0x18, 0x05, 0x20, 0x0E, 0x31, 0x1E, 0x2C, 0x3A,
	0x3B, 0x07, 0x58, 0x07, 0x1A, 0x00, 0x1B, 0x39, 0x01, 0x2B, 0x55, 0x13,
	0x0D, 0x39, 0x28, 0x2F, 0x51, 0x04, 0x2D, 0x7B, 0x01, 0x59, 0x1A, 0x5B,
	0x38, 0x1E, 0x57, 0x1B, 0x58, 0x13, 0x36, 0x0F, 0x2B, 0x04, 0x14, 0x22,
	0x0D, 0x37, 0x05, 0x06, 0x14, 0x11, 0x07, 0x05, 0x06, 0x35, 0x32, 0x1E,
	0x1A, 0x07, 0x5F, 0x37, 0x37, 0x3D, 0x72, 0x5E, 0x00, 0x18, 0x52, 0x11,
	0x59, 0x24, 0x37, 0x38, 0x0D, 0x34, 0x23, 0x26, 0x5B, 0x08, 0x29, 0x0C,
	0x5A, 0x22, 0x73, 0x06, 0x50, 0x06, 0x24, 0x75, 0x5F, 0x08, 0x2A, 0x21,
	0x14, 0x0D, 0x56, 0x29, 0x19, 0x36, 0x0D, 0x3B, 0x3E, 0x40, 0x25, 0x34,
	0x55, 0x23, 0x3E, 0x32, 0x06, 0x0F, 0x24, 0x18, 0x08, 0x24, 0x06, 0x29,
	0x2C, 0x35, 0x01, 0x14, 0x3F, 0x2F, 0x0C, 0x1D, 0x2B, 0x41, 0x11, 0x76,
	0x23, 0x0B, 0x59, 0x40, 0x08, 0x39, 0x57, 0x41, 0x27, 0x16, 0x01, 0x28,
	0x24, 0x5C, 0x3B, 0x15, 0x07, 0x34, 0x20, 0x11, 0x47, 0x07, 0x37, 0x1A,
	0x14, 0x2A, 0x0C, 0x3E, 0x19, 0x13, 0x43, 0x07, 0x04, 0x1B, 0x06, 0x59,
	0x56, 0x29, 0x07, 0x13, 0x1F, 0x2D, 0x5C, 0x24, 0x36, 0x28, 0x24, 0x5C,
	0x0E, 0x13, 0x21, 0x56, 0x21, 0x38, 0x05, 0x5B, 0x51, 0x59, 0x27, 0x0B,
	0x54, 0x38, 0x5C, 0x03, 0x12, 0x06, 0x03, 0x22, 0x11, 0x7A, 0x27, 0x02,
	0x1D, 0x58, 0x01, 0x1A, 0x33, 0x26, 0x0A, 0x29, 0x1C, 0x37, 0x1A, 0x44,
	0x13, 0x03, 0x32, 0x03, 0x3B, 0x38, 0x36, 0x54, 0x2D, 0x53, 0x17, 0x14,
	0x2A, 0x08, 0x58, 0x16, 0x0E, 0x28, 0x01, 0x2F, 0x75, 0x26, 0x2C, 0x3A,
	0x2D, 0x27, 0x0B, 0x0D, 0x28, 0x0F, 0x3B, 0x16, 0x14, 0x1E, 0x29, 0x74,
	0x5A, 0x53, 0x1E, 0x26, 0x07, 0x24, 0x24, 0x41, 0x59, 0x2E, 0x5D, 0x2D,
	0x45, 0x05, 0x10, 0x20, 0x06, 0x1B, 0x29, 0x27, 0x03, 0x2A, 0x20, 0x0D,
	0x2D, 0x28, 0x07, 0x1B, 0x31, 0x0C, 0x5B, 0x2B, 0x02, 0x0C, 0x16, 0x15,
	0x14, 0x22, 0x3F, 0x13, 0x5D, 0x0E, 0x23, 0x03, 0x38, 0x3D, 0x3B, 0x0A,
	0x21, 0x09, 0x5A, 0x08, 0x3C, 0x24, 0x69, 0x35, 0x27, 0x02, 0x1D, 0x05,
	0x2F, 0x05, 0x29, 0x07, 0x08, 0x0B, 0x04, 0x14, 0x2C, 0x0C, 0x5A, 0x08,
	0x21, 0x09, 0x37, 0x36, 0x58, 0x3E, 0x2E, 0x31, 0x1F, 0x25, 0x21, 0x38,
	0x10, 0x0F, 0x14, 0x08, 0x3E, 0x75, 0x1D, 0x09, 0x36, 0x3F, 0x0A, 0x5B,
	0x2C, 0x06, 0x27, 0x1B, 0x0D, 0x0B, 0x27, 0x2C, 0x1B, 0x1F, 0x58, 0x0F,
	0x3F, 0x01, 0x39, 0x14, 0x2F, 0x52, 0x36, 0x3B, 0x32, 0x24, 0x05, 0x04,
	0x03, 0x34, 0x3D, 0x23, 0x21, 0x19, 0x37, 0x3F, 0x09, 0x34, 0x25, 0x10,
	0x2B, 0x3D, 0x30, 0x3C, 0x27, 0x5F, 0x20, 0x74, 0x05, 0x2B, 0x0C, 0x0D,
	0x2A, 0x2A, 0x0F, 0x18, 0x32, 0x16, 0x00, 0x28, 0x17, 0x2E, 0x17, 0x34,
	0x04, 0x1C, 0x04, 0x29, 0x38, 0x51, 0x18, 0x27, 0x35, 0x07, 0x23, 0x06,
	0x5E, 0x05, 0x3C, 0x0D, 0x07, 0x3D, 0x11, 0x05, 0x26, 0x21, 0x0E, 0x31,
	0x02, 0x22, 0x1B, 0x00, 0x37, 0x2E, 0x23, 0x3D, 0x00, 0x37, 0x34, 0x39,
	0x25, 0x33, 0x34, 0x18, 0x0D, 0x02, 0x53, 0x2C, 0x43, 0x18, 0x0C, 0x21,
	0x7B, 0x34, 0x03, 0x5B, 0x25, 0x74, 0x19, 0x30, 0x05, 0x00, 0x00, 0x07,
	0x2D, 0x1E, 0x0E, 0x77, 0x08, 0x0F, 0x0D, 0x3D, 0x6D, 0x0E, 0x12, 0x20,
	0x5D, 0x06, 0x2D, 0x3B, 0x2C, 0x06, 0x32, 0x29, 0x29, 0x0F, 0x23, 0x01,
	0x38, 0x38, 0x02, 0x3A, 0x16, 0x00, 0x2B, 0x29, 0x31, 0x0C, 0x02, 0x0D,
	0x06, 0x04, 0x05, 0x25, 0x24, 0x5F, 0x09, 0x1A, 0x20, 0x0E, 0x2B, 0x2D,
	0x2D, 0x14, 0x0E, 0x25, 0x03, 0x15, 0x39, 0x26, 0x5E, 0x38, 0x74, 0x34,
	0x53, 0x0C, 0x1E, 0x36, 0x29, 0x1B, 0x17, 0x19, 0x07, 0x55, 0x23, 0x20,
	0x19, 0x24, 0x2B, 0x00, 0x59, 0x19, 0x23, 0x5A, 0x39, 0x36, 0x02, 0x72,
	0x24, 0x15, 0x34, 0x33, 0x7A, 0x04, 0x03, 0x01, 0x53, 0x7B, 0x2A, 0x50,
	0x5B, 0x20, 0x2E, 0x05, 0x25, 0x04, 0x5D, 0x3A, 0x3B, 0x54, 0x38, 0x25,
	0x2A, 0x1C, 0x3B, 0x26, 0x1B, 0x04, 0x21, 0x38, 0x26, 0x0E, 0x0A, 0x58,
	0x25, 0x0D, 0x01, 0x15, 0x1A, 0x36, 0x3E, 0x3F, 0x29, 0x1F, 0x37, 0x06,
	0x19, 0x7B, 0x27, 0x00, 0x2D, 0x09, 0x0D, 0x2B, 0x34, 0x18, 0x0E, 0x2F,
	0x47, 0x38, 0x21, 0x31, 0x16, 0x0E, 0x0E, 0x39, 0x3C, 0x1B, 0x35, 0x11,
	0x2C, 0x22, 0x7B, 0x2F, 0x2F, 0x2C, 0x59, 0x17, 0x20, 0x14, 0x3D, 0x59,
	0x13, 0x1D, 0x0A, 0x08, 0x26, 0x07, 0x20, 0x2B, 0x29, 0x23, 0x2D, 0x2D,
	0x39, 0x39, 0x13, 0x0D, 0x26, 0x34, 0x26, 0x3B, 0x21, 0x0A, 0x0A, 0x34,
	0x0D, 0x12, 0x23, 0x06, 0x5A, 0x06, 0x0C, 0x16, 0x29, 0x3B, 0x12, 0x15,
	0x59, 0x2B, 0x2C, 0x0F, 0x71, 0x1D, 0x52, 0x3C, 0x0C, 0x16, 0x5F, 0x0B,
	0x03, 0x27, 0x73, 0x0E, 0x10, 0x17, 0x2A, 0x20, 0x5A, 0x29, 0x2C, 0x01,
	0x2D, 0x5D, 0x08, 0x17, 0x2C, 0x2E, 0x29, 0x13, 0x3A, 0x1F, 0x1A, 0x3A,
	0x4E, 0x29, 0x07, 0x0A, 0x29, 0x26, 0x5B, 0x32, 0x71, 0x15, 0x00, 0x2A,
	0x2E, 0x20, 0x06, 0x4E, 0x1A, 0x24, 0x00, 0x09, 0x30, 0x3B, 0x22, 0x24,
	0x3D, 0x28, 0x5F, 0x5D, 0x2E, 0x5A, 0x05, 0x5B, 0x0A, 0x32, 0x27, 0x0E,
	0x0F, 0x12, 0x18, 0x58, 0x04, 0x5B, 0x1A, 0x24, 0x43, 0x06, 0x20, 0x0C,
	0x06, 0x39, 0x20, 0x39, 0x31, 0x31, 0x43, 0x22, 0x3A, 0x0C, 0x06, 0x3D,
	0x51, 0x41, 0x2E, 0x0F, 0x1E, 0x18, 0x25, 0x07, 0x32, 0x08, 0x17, 0x02,
	0x09, 0x18, 0x5D, 0x23, 0x0B, 0x13, 0x73, 0x2E, 0x4A, 0x14, 0x1D, 0x7B,
	0x1A, 0x55, 0x25, 0x59, 0x08, 0x2A, 0x05, 0x25, 0x58, 0x16, 0x35, 0x2D,
	0x00, 0x02, 0x6D, 0x5D, 0x4E, 0x19, 0x13, 0x36, 0x55, 0x52, 0x5C, 0x2E,
	0x32, 0x06, 0x20, 0x1D, 0x23, 0x13, 0x2E, 0x09, 0x22, 0x3B, 0x2E, 0x16,
	0x11, 0x1B, 0x2D, 0x37, 0x59, 0x14, 0x5B, 0x2A, 0x09, 0x2A, 0x03, 0x3E,
	0x29, 0x35, 0x3C, 0x14, 0x0D, 0x28, 0x08, 0x2F, 0x17, 0x56, 0x05, 0x2F,
	0x23, 0x17, 0x27, 0x2A, 0x0D, 0x39, 0x2E, 0x56, 0x0E, 0x15, 0x1F, 0x10,
	0x57, 0x0E, 0x3A, 0x03, 0x3B, 0x5A, 0x24, 0x30, 0x0F, 0x03, 0x07, 0x00,
	0x0F, 0x29, 0x0E, 0x25, 0x1D, 0x14, 0x1D, 0x54, 0x09, 0x2A, 0x25, 0x27,
	0x39, 0x3B, 0x2A, 0x70, 0x19, 0x32, 0x17, 0x1C, 0x0E, 0x22, 0x0E, 0x21,
	0x25, 0x03, 0x1A, 0x11, 0x09, 0x32, 0x7A, 0x06, 0x07, 0x07, 0x05, 0x31,
	0x2F, 0x54, 0x2B, 0x12, 0x04, 0x5F, 0x17, 0x2F, 0x40, 0x17, 0x22, 0x53,
	0x5B, 0x58, 0x12, 0x3C, 0x51, 0x04, 0x2A, 0x0C, 0x2F, 0x14, 0x22, 0x08,
	0x2D, 0x08, 0x14, 0x41, 0x06, 0x0A, 0x19, 0x54, 0x5F, 0x2C, 0x70, 0x55,
	0x55, 0x21, 0x00, 0x0A, 0x14, 0x03, 0x56, 0x3B, 0x16, 0x5D, 0x50, 0x2B,
	0x59, 0x1B, 0x3A, 0x52, 0x21, 0x2F, 0x16, 0x29, 0x28, 0x0A, 0x04, 0x77,
	0x21, 0x38, 0x06, 0x59, 0x10, 0x14, 0x0B, 0x3C, 0x3A, 0x12, 0x24, 0x23,
	0x07, 0x0F, 0x31, 0x3E, 0x51, 0x0F, 0x3A, 0x0B, 0x03, 0x11, 0x5E, 0x00,
	0x3B, 0x3C, 0x2E, 0x2A, 0x27, 0x3B, 0x35, 0x27, 0x58, 0x21, 0x73, 0x27,
	0x50, 0x2D, 0x44, 0x24, 0x1D, 0x0C, 0x2F, 0x3C, 0x74, 0x05, 0x33, 0x2A,
	0x29, 0x0F, 0x5D, 0x06, 0x08, 0x19, 0x28, 0x1C, 0x0A, 0x03, 0x40, 0x16,
	0x5B, 0x51, 0x1E, 0x27, 0x10, 0x2F, 0x28, 0x3E, 0x19, 0x07, 0x3F, 0x03,
	0x1E, 0x5C, 0x13, 0x16, 0x05, 0x24, 0x5C, 0x26, 0x5D, 0x06, 0x29, 0x0F,
	0x32, 0x14, 0x2E, 0x3A, 0x26, 0x2E, 0x3A, 0x0A, 0x2B, 0x29, 0x77, 0x0A,
	0x08, 0x0C, 0x59, 0x1B, 0x0F, 0x08, 0x1F, 0x32, 0x31, 0x1A, 0x05, 0x0C,
	0x3A, 0x29, 0x1B, 0x17, 0x08, 0x32, 0x00, 0x5B, 0x27, 0x25, 0x3A, 0x2E,
	0x2E, 0x0A, 0x0F, 0x59, 0x0F, 0x38, 0x50, 0x27, 0x3D, 0x00, 0x27, 0x0E,
	0x14, 0x3C, 0x05, 0x58, 0x06, 0x5B, 0x26, 0x00, 0x07, 0x2B, 0x16, 0x5B,
	0x12, 0x28, 0x25, 0x01, 0x2F, 0x0D, 0x0D, 0x27, 0x41, 0x3F, 0x70, 0x58,
	0x05, 0x3D, 0x31, 0x34, 0x2E, 0x38, 0x37, 0x3A, 0x0D, 0x24, 0x20, 0x25,
	0x1F, 0x23, 0x23, 0x07, 0x59, 0x0D, 0x0E, 0x3A, 0x36, 0x07, 0x26, 0x2C,
	0x38, 0x0A, 0x36, 0x3C, 0x00, 0x55, 0x2A, 0x2A, 0x5C, 0x70, 0x22, 0x59,
	0x18, 0x0F, 0x3B, 0x0B, 0x11, 0x1E, 0x52, 0x29, 0x09, 0x52, 0x14, 0x00,
	0x75, 0x2D, 0x2F, 0x0B, 0x2D, 0x7B, 0x0B, 0x02, 0x22, 0x0F, 0x21, 0x54,
	0x0E, 0x1F, 0x52, 0x18, 0x0F, 0x29, 0x57, 0x21, 0x71, 0x1C, 0x09, 0x00,
	0x00, 0x2C, 0x29, 0x52, 0x25, 0x0E, 0x0D, 0x07, 0x00, 0x2F, 0x2D, 0x31,
	0x1B, 0x0F, 0x05, 0x3A, 0x3A, 0x01, 0x39, 0x59, 0x2A, 0x2A, 0x09, 0x05,
	0x04, 0x18, 0x20, 0x5D, 0x55, 0x26, 0x5C, 0x16, 0x34, 0x36, 0x03, 0x5E,
	0x23, 0x00, 0x51, 0x22, 0x59, 0x2A, 0x2A, 0x55, 0x41, 0x18, 0x30, 0x06,
	0x06, 0x56, 0x32, 0x04, 0x38, 0x1B, 0x0C, 0x1E, 0x09, 0x39, 0x51, 0x59,
	0x04, 0x69, 0x29, 0x25, 0x1A, 0x0E, 0x34, 0x59, 0x08, 0x29, 0x19, 0x76,
	0x39, 0x2D, 0x45, 0x33, 0x26, 0x2A, 0x36, 0x09, 0x1D, 0x0C, 0x15, 0x58,
	0x3C, 0x18, 0x69, 0x2E, 0x30, 0x20, 0x29, 0x14, 0x5F, 0x38, 0x14, 0x18,
	0x71, 0x19, 0x2C, 0x09, 0x23, 0x77, 0x59, 0x54, 0x2A, 0x3D, 0x0C, 0x15,
	0x27, 0x16, 0x28, 0x75, 0x1E, 0x0C, 0x0D, 0x12, 0x13, 0x5C, 0x02, 0x17,
	0x3A, 0x71, 0x2E, 0x07, 0x08, 0x2A, 0x1B, 0x26, 0x15, 0x05, 0x23, 0x7B,
	0x55, 0x06, 0x3F, 0x5B, 0x2C, 0x14, 0x10, 0x16, 0x24, 0x69, 0x22, 0x00,
	0x59, 0x39, 0x30, 0x0E, 0x10, 0x00, 0x25, 0x31, 0x0B, 0x36, 0x22, 0x0A,
	0x37, 0x2E, 0x0E, 0x5B, 0x29, 0x35, 0x28, 0x03, 0x1C, 0x40, 0x37, 0x07,
	0x1B, 0x0D, 0x59, 0x36, 0x1E, 0x2C, 0x5F, 0x5C, 0x31, 0x0F, 0x51, 0x17,
	0x0D, 0x0F, 0x24, 0x25, 0x0D, 0x2F, 0x2A, 0x5F, 0x31, 0x56, 0x5A, 0x26,
	0x24, 0x54, 0x5A, 0x5C, 0x21, 0x28, 0x14, 0x37, 0x44, 0x2F, 0x19, 0x55,
	0x5A, 0x5E, 0x20, 0x04, 0x33, 0x41, 0x09, 0x08, 0x25, 0x0C, 0x23, 0x11,
	0x09, 0x07, 0x0C, 0x20, 0x0A, 0x29, 0x3D, 0x50, 0x07, 0x0C, 0x76, 0x5A,
	0x2F, 0x3D, 0x32, 0x07, 0x29, 0x0A, 0x58, 0x39, 0x0D, 0x06, 0x33, 0x1A,
	0x25, 0x1B, 0x35, 0x39, 0x06, 0x0E, 0x24, 0x5F, 0x31, 0x0C, 0x1B, 0x3B,
	0x00, 0x03, 0x14, 0x03, 0x0C, 0x26, 0x10, 0x3F, 0x5F, 0x0E, 0x07, 0x59,
	0x23, 0x1B, 0x30, 0x03, 0x38, 0x2B, 0x31, 0x03, 0x43, 0x55, 0x2B, 0x05,
	0x35, 0x02, 0x0E, 0x14, 0x26, 0x2A, 0x5B, 0x33, 0x5F, 0x0F, 0x18, 0x3A,
	0x04, 0x3E, 0x5E, 0x0C, 0x55, 0x23, 0x57, 0x5D, 0x06, 0x36, 0x02, 0x26,
	0x3B, 0x33, 0x24, 0x0D, 0x21, 0x5D, 0x30, 0x09, 0x05, 0x17, 0x20, 0x74,
	0x06, 0x25, 0x5B, 0x08, 0x3A, 0x0B, 0x29, 0x19, 0x03, 0x74, 0x5F, 0x07,
	0x07, 0x5F, 0x10, 0x19, 0x0E, 0x5A, 0x29, 0x2E, 0x22, 0x05, 0x05, 0x12,
	0x33, 0x05, 0x30, 0x22, 0x22, 0x0C, 0x2E, 0x11, 0x3F, 0x03, 0x1B, 0x1C,
	0x2D, 0x3A, 0x44, 0x20, 0x3E, 0x50, 0x23, 0x21, 0x30, 0x25, 0x07, 0x3D,
	0x0F, 0x34, 0x02, 0x0F, 0x19, 0x26, 0x03, 0x16, 0x53, 0x03, 0x12, 0x70,
	0x04, 0x36, 0x0A, 0x3F, 0x73, 0x02, 0x24, 0x5C, 0x23, 0x75, 0x20, 0x3B,
	0x08, 0x2D, 0x29, 0x09, 0x2E, 0x5B, 0x18, 0x03, 0x16, 0x38, 0x34, 0x44,
	0x33, 0x00, 0x1B, 0x04, 0x12, 0x2B, 0x1E, 0x39, 0x0D, 0x3F, 0x20, 0x3C,
	0x30, 0x1D, 0x3C, 0x03, 0x3E, 0x24, 0x19, 0x59, 0x18, 0x03, 0x24, 0x03,
	0x07, 0x31, 0x0F, 0x14, 0x3B, 0x21, 0x77, 0x05, 0x18, 0x07, 0x13, 0x2C,
	0x18, 0x26, 0x2A, 0x38, 0x23, 0x39, 0x28, 0x5D, 0x0F, 0x2C, 0x00, 0x12,
	0x1E, 0x52, 0x2B, 0x29, 0x07, 0x36, 0x52, 0x01, 0x3B, 0x50, 0x0B, 0x0D,
	0x1B, 0x01, 0x15, 0x38, 0x33, 0x03, 0x39, 0x17, 0x34, 0x5E, 0x69, 0x07,
	0x12, 0x37, 0x18, 0x18, 0x2A, 0x3B, 0x1F, 0x0E, 0x3B, 0x1B, 0x3B, 0x21,
	0x25, 0x00, 0x29, 0x1B, 0x45, 0x00, 0x23, 0x1F, 0x55, 0x45, 0x3C, 0x20,
	0x15, 0x10, 0x06, 0x33, 0x16, 0x04, 0x17, 0x45, 0x32, 0x16, 0x3F, 0x28,
	0x04, 0x0F, 0x7B, 0x2F, 0x28, 0x06, 0x2A, 0x71, 0x58, 0x15, 0x18, 0x23,
	0x1A, 0x29, 0x1B, 0x00, 0x05, 0x0C, 0x36, 0x54, 0x00, 0x3A, 0x20, 0x18,
	0x0A, 0x0A, 0x03, 0x77, 0x14, 0x02, 0x05, 0x04, 0x34, 0x06, 0x36, 0x01,
	0x3F, 0x18, 0x3B, 0x30, 0x57, 0x2C, 0x1B, 0x1E, 0x0C, 0x1A, 0x3D, 0x71,
	0x00, 0x54, 0x20, 0x31, 0x24, 0x3D, 0x17, 0x0B, 0x58, 0x76, 0x39, 0x09,
	0x3F, 0x0E, 0x2D, 0x28, 0x25, 0x39, 0x12, 0x6D, 0x3B, 0x06, 0x17, 0x26,
	0x12, 0x35, 0x0A, 0x28, 0x19, 0x2F, 0x35, 0x27, 0x0D, 0x19, 0x13, 0x2F,
	0x4A, 0x36, 0x01, 0x0F, 0x21, 0x37, 0x0B, 0x52, 0x10, 0x05, 0x14, 0x38,
	0x3F, 0x77, 0x3D, 0x35, 0x0F, 0x2F, 0x74, 0x2A, 0x33, 0x36, 0x1E, 0x3A,
	0x03, 0x15, 0x5C, 0x03, 0x33, 0x26, 0x0E, 0x25, 0x29, 0x13, 0x26, 0x31,
	0x0F, 0x44, 0x0D, 0x0A, 0x08, 0x08, 0x5A, 0x26, 0x5F, 0x02, 0x1E, 0x0E,
	0x2B, 0x1A, 0x29, 0x02, 0x02, 0x32, 0x3C, 0x15, 0x20, 0x1A, 0x3B, 0x58,
	0x57, 0x20, 0x5D, 0x36, 0x35, 0x10, 0x01, 0x1E, 0x35, 0x54, 0x55, 0x5C,
	0x1E, 0x14, 0x1C, 0x54, 0x37, 0x0D, 0x20, 0x59, 0x56, 0x2A, 0x38, 0x73,
	0x1D, 0x32, 0x41, 0x04, 0x74, 0x18, 0x39, 0x07, 0x44, 0x1B, 0x35, 0x32,
	0x3B, 0x3D, 0x21, 0x3A, 0x00, 0x02, 0x38, 0x0F, 0x3F, 0x59, 0x01, 0x32,
	0x30, 0x36, 0x53, 0x1A, 0x1C, 0x72, 0x5F, 0x23, 0x20, 0x40, 0x07, 0x22,
	0x13, 0x0A, 0x27, 0x1B, 0x54, 0x52, 0x3E, 0x39, 0x12, 0x38, 0x36, 0x5E,
	0x28, 0x35, 0x1D, 0x16, 0x3A, 0x08, 0x14, 0x35, 0x08, 0x2F, 0x52, 0x34,
	0x5F, 0x13, 0x1A, 0x40, 0x27, 0x2B, 0x33, 0x07, 0x06, 0x00, 0x39, 0x57,
	0x3A, 0x59, 0x20, 0x18, 0x11, 0x3B, 0x31, 0x37, 0x20, 0x16, 0x1D, 0x19,
	0x18, 0x0D, 0x00, 0x0B, 0x31, 0x1A, 0x1E, 0x00, 0x3C, 0x12, 0x30, 0x28,
	0x00, 0x2A, 0x40, 0x35, 0x24, 0x39, 0x36, 0x3D, 0x74, 0x05, 0x39, 0x20,
	0x2D, 0x12, 0x1C, 0x12, 0x09, 0x20, 0x16, 0x0B, 0x23, 0x5F, 0x2F, 0x29,
	0x3D, 0x15, 0x0C, 0x0C, 0x1A, 0x06, 0x59, 0x5F, 0x0A, 0x12, 0x08, 0x0B,
	0x2C, 0x0E, 0x0C, 0x47, 0x31, 0x56, 0x33, 0x04, 0x07, 0x1B, 0x2D, 0x02,
	0x25, 0x20, 0x34, 0x1F, 0x2C, 0x75, 0x35, 0x4E, 0x2C, 0x3D, 0x17, 0x07,
	0x0A, 0x2C, 0x12, 0x11, 0x5D, 0x58, 0x2D, 0x27, 0x1B, 0x1A, 0x1B, 0x39,
	0x1A, 0x28, 0x1A, 0x4A, 0x1E, 0x24, 0x23, 0x47, 0x06, 0x19, 0x1A, 0x00,
	0x21, 0x32, 0x3A, 0x01, 0x28, 0x26, 0x58, 0x07, 0x31, 0x21, 0x34, 0x51,
	0x23, 0x01, 0x76, 0x1F, 0x2F, 0x37, 0x27, 0x30, 0x5E, 0x33, 0x2D, 0x03,
	0x23, 0x35, 0x34, 0x08, 0x25, 0x21, 0x0E, 0x0D, 0x08, 0x06, 0x18, 0x5D,
	0x24, 0x56, 0x20, 0x0D, 0x5A, 0x57, 0x22, 0x2D, 0x2E, 0x0B, 0x03, 0x21,
	0x32, 0x1A, 0x1F, 0x3B, 0x5C, 0x53, 0x7A, 0x2E, 0x0C, 0x2A, 0x40, 0x7A,
	0x2B, 0x0E, 0x5C, 0x33, 0x16, 0x59, 0x00, 0x2A, 0x53, 0x26, 0x26, 0x26,
	0x3F, 0x38, 0x0A, 0x2B, 0x36, 0x58, 0x07, 0x04, 0x3C, 0x11, 0x57, 0x0A,
	0x7B, 0x2D, 0x14, 0x1B, 0x3E, 0x38, 0x16, 0x2E, 0x22, 0x05, 0x17, 0x54,
	0x17, 0x2F, 0x25, 0x35, 0x02, 0x00, 0x02, 0x5F, 0x00, 0x05, 0x2F, 0x28,
	0x26, 0x16, 0x5F, 0x06, 0x34, 0x5B, 0x2A, 0x1F, 0x56, 0x37, 0x21, 0x25,
	0x19, 0x23, 0x59, 0x0E, 0x06, 0x26, 0x1B, 0x03, 0x00, 0x21, 0x55, 0x1B,
	0x45, 0x2F, 0x32, 0x58, 0x13, 0x07, 0x1F, 0x28, 0x5B, 0x02, 0x08, 0x11,
	0x2D, 0x26, 0x15, 0x2B, 0x1A, 0x03, 0x29, 0x0C, 0x41, 0x09, 0x6D, 0x1B,
	0x0F, 0x2F, 0x12, 0x37, 0x2A, 0x0A, 0x18, 0x24, 0x29, 0x22, 0x0F, 0x19,
	0x44, 0x05, 0x5B, 0x0E, 0x01, 0x5C, 0x29, 0x3D, 0x30, 0x5D, 0x09, 0x33,
	0x3B, 0x03, 0x07, 0x01, 0x01, 0x2D, 0x03, 0x5F, 0x44, 0x25, 0x2F, 0x2E,
	0x1B, 0x5A, 0x72, 0x58, 0x26, 0x3C, 0x5A, 0x21, 0x47, 0x16, 0x22, 0x2C,
	0x0B, 0x34, 0x06, 0x29, 0x1F, 0x23, 0x2A, 0x2B, 0x45, 0x39, 0x1A, 0x54,
	0x09, 0x00, 0x1B, 0x7B, 0x5E, 0x1B, 0x3C, 0x40, 0x31, 0x07, 0x13, 0x26,
	0x1E, 0x24, 0x20, 0x04, 0x06, 0x2E, 0x11, 0x47, 0x0A, 0x02, 0x44, 0x25,
	0x35, 0x55, 0x1D, 0x04, 0x37, 0x2A, 0x14, 0x2C, 0x3B, 0x73, 0x38, 0x18,
	0x23, 0x40, 0x07, 0x08, 0x22, 0x3D, 0x22, 0x13, 0x1C, 0x24, 0x2D, 0x26,
	0x38, 0x2D, 0x05, 0x56, 0x27, 0x09, 0x28, 0x0F, 0x26, 0x5D, 0x23, 0x39,
	0x55, 0x41, 0x1E, 0x20, 0x27, 0x33, 0x5E, 0x2A, 0x3A, 0x18, 0x1B, 0x00,
	0x0E, 0x38, 0x5C, 0x39, 0x29, 0x58, 0x0D, 0x3A, 0x37, 0x01, 0x5A, 0x31,
	0x5E, 0x17, 0x5E, 0x05, 0x16, 0x38, 0x2E, 0x5F, 0x40, 0x11, 0x0A, 0x00,
	0x5F, 0x09, 0x27, 0x3A, 0x0F, 0x29, 0x0A, 0x16, 0x24, 0x00, 0x01, 0x27,
	0x3A, 0x5E, 0x50, 0x37, 0x06, 0x35, 0x1A, 0x32, 0x0D, 0x25, 0x09, 0x58,
	0x17, 0x39, 0x2A, 0x0A, 0x58, 0x0B, 0x26, 0x09, 0x11, 0x00, 0x13, 0x3C,
	0x33, 0x11, 0x5C, 0x59, 0x3E, 0x1C, 0x36, 0x3F, 0x13, 0x18, 0x0F, 0x09,
	0x26, 0x09, 0x2C, 0x5E, 0x33, 0x01, 0x35, 0x34, 0x20, 0x0E, 0x04, 0x16,
	0x20, 0x12, 0x04, 0x01, 0x07, 0x58, 0x38, 0x7B, 0x2B, 0x37, 0x56, 0x31,
	0x37, 0x58, 0x26, 0x3F, 0x2E, 0x28, 0x16, 0x52, 0x1C, 0x44, 0x3A, 0x34,
	0x54, 0x3D, 0x13, 0x37, 0x01, 0x0A, 0x36, 0x07, 0x2A, 0x19, 0x50, 0x5D,
	0x1C, 0x23, 0x5F, 0x0E, 0x19, 0x02, 0x18, 0x1E, 0x2B, 0x28, 0x19, 0x11,
	0x34, 0x37, 0x03, 0x2D, 0x0C, 0x5E, 0x2E, 0x2D, 0x03, 0x11, 0x02, 0x2C,
	0x0B, 0x04, 0x35, 0x5E, 0x36, 0x2D, 0x06, 0x15, 0x28, 0x13, 0x07, 0x39,
	0x0A, 0x0D, 0x35, 0x24, 0x19, 0x09, 0x08, 0x33, 0x5C, 0x12, 0x72, 0x1C,
	0x16, 0x16, 0x05, 0x18, 0x3F, 0x0F, 0x0C, 0x01, 0x72, 0x07, 0x08, 0x58,
	0x33, 0x6D, 0x58, 0x04, 0x02, 0x1D, 0x7A, 0x5C, 0x2D, 0x01, 0x12, 0x31,
	0x2F, 0x12, 0x3D, 0x2F, 0x0F, 0x3D, 0x18, 0x14, 0x59, 0x20, 0x3B, 0x16,
	0x18, 0x28, 0x2D, 0x43, 0x23, 0x16, 0x59, 0x04, 0x0D, 0x51, 0x07, 0x3D,
	0x21, 0x2A, 0x2E, 0x01, 0x33, 0x2A, 0x02, 0x11, 0x38, 0x05, 0x7A, 0x22,
	0x08, 0x0C, 0x24, 0x06, 0x0A, 0x35, 0x1D, 0x5C, 0x12, 0x1B, 0x31, 0x5C,
	0x28, 0x69, 0x1F, 0x17, 0x1C, 0x19, 0x0D, 0x58, 0x27, 0x34, 0x0C, 0x7B,
	0x0B, 0x19, 0x2A, 0x1A, 0x6D, 0x16, 0x06, 0x08, 0x01, 0x12, 0x3D, 0x06,
	0x34, 0x12, 0x0F, 0x28, 0x05, 0x3C, 0x3C, 0x74, 0x2B, 0x2D, 0x2B, 0x13,
	0x03, 0x06, 0x32, 0x0F, 0x1A, 0x73, 0x5F, 0x16, 0x20, 0x03, 0x0F, 0x22,
	0x51, 0x29, 0x3C, 0x01, 0x5A, 0x56, 0x23, 0x59, 0x77, 0x1F, 0x4A, 0x38,
	0x2A, 0x77, 0x27, 0x59, 0x39, 0x52, 0x70, 0x5F, 0x29, 0x5E, 0x24, 0x11,
	0x21, 0x31, 0x37, 0x18, 0x28, 0x0B, 0x2D, 0x39, 0x02, 0x0A, 0x20, 0x0C,
	0x34, 0x11, 0x7A, 0x05, 0x23, 0x0F, 0x38, 0x26, 0x3D, 0x10, 0x34, 0x0C,
	0x6D, 0x23, 0x38, 0x26, 0x07, 0x04, 0x5D, 0x13, 0x2C, 0x0D, 0x27, 0x1C,
	0x51, 0x56, 0x03, 0x74, 0x28, 0x52, 0x57, 0x22, 0x0A, 0x03, 0x50, 0x02,
	0x32, 0x01, 0x05, 0x10, 0x26, 0x52, 0x13, 0x2E, 0x06, 0x57, 0x5A, 0x75,
	0x3B, 0x11, 0x3E, 0x2F, 0x25, 0x3C, 0x2B, 0x3E, 0x44, 0x17, 0x05, 0x03,
	0x24, 0x0D, 0x6D, 0x59, 0x59, 0x0F, 0x53, 0x3A, 0x34, 0x55, 0x20, 0x0F,
	0x34, 0x5A, 0x22, 0x5B, 0x3A, 0x71, 0x1B, 0x29, 0x03, 0x5A, 0x7A, 0x05,
	0x16, 0x37, 0x44, 0x05, 0x09, 0x00, 0x2A, 0x3F, 0x7B, 0x36, 0x0E, 0x56,
	0x0C, 0x15, 0x2B, 0x53, 0x56, 0x59, 0x75, 0x1E, 0x1B, 0x29, 0x07, 0x32,
	0x27, 0x39, 0x01, 0x3C, 0x74, 0x08, 0x52, 0x5B, 0x3D, 0x12, 0x59, 0x14,
	0x2A, 0x22, 0x77, 0x1B, 0x17, 0x27, 0x0A, 0x2E, 0x5F, 0x17, 0x28, 0x20,
	0x6D, 0x2F, 0x22, 0x0D, 0x1C, 0x15, 0x2D, 0x2B, 0x21, 0x01, 0x01, 0x3C,
	0x04, 0x1F, 0x22, 0x76, 0x21, 0x37, 0x59, 0x23, 0x23, 0x3B, 0x25, 0x57,
	0x12, 0x72, 0x01, 0x27, 0x14, 0x58, 0x0A, 0x54, 0x26, 0x5D, 0x1C, 0x0B,
	0x28, 0x2A, 0x0D, 0x32, 0x04, 0x2A, 0x10, 0x25, 0x24, 0x6D, 0x0E, 0x58,
	0x5B, 0x3D, 0x09, 0x0F, 0x4E, 0x19, 0x26, 0x37, 0x14, 0x33, 0x1D, 0x0C,
	0x3A, 0x2D, 0x2D, 0x3E, 0x05, 0x36, 0x20, 0x51, 0x36, 0x0A, 0x6D, 0x14,
	0x16, 0x1A, 0x5F, 0x03, 0x43, 0x03, 0x5C, 0x19, 0x29, 0x2D, 0x0D, 0x08,
	0x53, 0x01, 0x5C, 0x16, 0x5A, 0x3F, 0x7B, 0x25, 0x4E, 0x2A, 0x3C, 0x2D,
	0x3A, 0x06, 0x57, 0x11, 0x2A, 0x29, 0x04, 0x21, 0x12, 0x12, 0x5F, 0x27,
	0x0B, 0x2C, 0x12, 0x35, 0x1B, 0x57, 0x27, 0x34, 0x43, 0x54, 0x0F, 0x01,
	0x3A, 0x1F, 0x38, 0x0B, 0x02, 0x0F, 0x1C, 0x30, 0x18, 0x2F, 0x0C, 0x26,
	0x4E, 0x3C, 0x11, 0x26, 0x3B, 0x2C, 0x1F, 0x5A, 0x2C, 0x0E, 0x25, 0x21,
	0x1B, 0x74, 0x2F, 0x19, 0x19, 0x2E, 0x04, 0x3F, 0x02, 0x41, 0x05, 0x0A,
	0x1A, 0x57, 0x0B, 0x5F, 0x27, 0x15, 0x03, 0x3B, 0x0D, 0x0D, 0x03, 0x15,
	0x3C, 0x5B, 0x25, 0x27, 0x39, 0x37, 0x04, 0x2E, 0x5D, 0x13, 0x36, 0x3A,
	0x38, 0x1A, 0x0D, 0x01, 0x27, 0x0D, 0x2A, 0x2F, 0x5A, 0x1F, 0x11, 0x3A,
	0x16, 0x27, 0x18, 0x06, 0x1E, 0x57, 0x2B, 0x3C, 0x17, 0x0F, 0x0D, 0x08,
	0x44, 0x06, 0x5E, 0x35, 0x3E, 0x04, 0x05, 0x59, 0x13, 0x08, 0x3F, 0x27,
	0x20, 0x4E, 0x14, 0x40, 0x04, 0x24, 0x0D, 0x2C, 0x04, 0x0B, 0x07, 0x0A,
	0x0C, 0x24, 0x0B, 0x47, 0x2E, 0x1A, 0x27, 0x0F, 0x26, 0x55, 0x0F, 0x09,
	0x2F, 0x29, 0x2D, 0x1D, 0x3B, 0x0E, 0x3A, 0x11, 0x24, 0x0E, 0x10, 0x55,
	0x26, 0x2D, 0x44, 0x3B, 0x0F, 0x39, 0x56, 0x52, 0x75, 0x2F, 0x31, 0x3C,
	0x3A, 0x32, 0x35, 0x37, 0x08, 0x1D, 0x31, 0x27, 0x24, 0x26, 0x3C, 0x04,
	0x2F, 0x1B, 0x2F, 0x0D, 0x3A, 0x3A, 0x1B, 0x36, 0x58, 0x2F, 0x38, 0x08,
	0x18, 0x3B, 0x07, 0x08, 0x03, 0x38, 0x09, 0x12, 0x5A, 0x22, 0x1C, 0x1A,
	0x69, 0x3C, 0x0F, 0x04, 0x53, 0x10, 0x1D, 0x0D, 0x18, 0x29, 0x24, 0x0B,
	0x20, 0x0D, 0x25, 0x76, 0x55, 0x13, 0x1B, 0x1C, 0x17, 0x2D, 0x32, 0x0A,
	0x1F, 0x0E, 0x0B, 0x31, 0x36, 0x0C, 0x23, 0x3E, 0x34, 0x41, 0x1C, 0x26,
	0x39, 0x0A, 0x0F, 0x11, 0x76, 0x2E, 0x57, 0x2F, 0x29, 0x32, 0x20, 0x39,
	0x0A, 0x23, 0x29, 0x3D, 0x4E, 0x3D, 0x1D, 0x05, 0x20, 0x57, 0x2C, 0x1B,
	0x09, 0x59, 0x0D, 0x08, 0x00, 0x34, 0x09, 0x0C, 0x56, 0x0A, 0x08, 0x0F,
	0x58, 0x5F, 0x25, 0x2B, 0x02, 0x2D, 0x5A, 0x2A, 0x7B, 0x03, 0x10, 0x05,
	0x2C, 0x0A, 0x25, 0x11, 0x0F, 0x02, 0x13, 0x2A, 0x04, 0x3A, 0x25, 0x1B,
	0x05, 0x08, 0x38, 0x5C, 0x2B, 0x0F, 0x0F, 0x24, 0x1E, 0x69, 0x16, 0x18,
	0x18, 0x05, 0x1B, 0x09, 0x2F, 0x26, 0x40, 0x31, 0x2E, 0x18, 0x5F, 0x0F,
	0x14, 0x24, 0x28, 0x23, 0x20, 0x6D, 0x54, 0x11, 0x3E, 0x1A, 0x2D, 0x2F,
	0x1B, 0x5B, 0x00, 0x27, 0x38, 0x2D, 0x25, 0x3C, 0x75, 0x2B, 0x34, 0x0B,
	0x1F, 0x09, 0x2B, 0x2F, 0x3F, 0x3C, 0x0D, 0x5C, 0x31, 0x26, 0x3A, 0x00,
	0x01, 0x10, 0x0F, 0x3E, 0x2D, 0x3B, 0x2A, 0x3B, 0x0C, 0x2E, 0x54, 0x50,
	0x3F, 0x25, 0x0A, 0x19, 0x12, 0x18, 0x52, 0x74, 0x14, 0x03, 0x2B, 0x44,
	0x2C, 0x14, 0x52, 0x03, 0x1A, 0x3B, 0x04, 0x2A, 0x3C, 0x04, 0x37, 0x0F,
	0x0B, 0x18, 0x27, 0x36, 0x16, 0x19, 0x0A, 0x0F, 0x73, 0x47, 0x03, 0x1F,
	0x5C, 0x03, 0x03, 0x05, 0x06, 0x33, 0x72, 0x1F, 0x2E, 0x02, 0x0A, 0x75,
	0x36, 0x3B, 0x41, 0x01, 0x0D, 0x14, 0x0B, 0x19, 0x58, 0x76, 0x5F, 0x53,
	0x2F, 0x03, 0x28, 0x18, 0x2D, 0x3D, 0x18, 0x74, 0x02, 0x25, 0x21, 0x26,
	0x0A, 0x3F, 0x05, 0x1C, 0x22, 0x1A, 0x27, 0x4A, 0x0F, 0x3C, 0x2A, 0x3A,
	0x55, 0x21, 0x5D, 0x35, 0x34, 0x08, 0x45, 0x5D, 0x09, 0x04, 0x31, 0x28,
	0x00, 0x2A, 0x28, 0x14, 0x08, 0x1C, 0x37, 0x09, 0x32, 0x03, 0x38, 0x1B,
	0x1E, 0x0F, 0x25, 0x11, 0x38, 0x0E, 0x2B, 0x20, 0x53, 0x0A, 0x15, 0x2E,
	0x29, 0x13, 0x06, 0x2F, 0x24, 0x38, 0x40, 0x70, 0x38, 0x4A, 0x04, 0x2D,
	0x75, 0x5D, 0x14, 0x21, 0x3B, 0x05, 0x08, 0x34, 0x27, 0x07, 0x76, 0x27,
	0x0A, 0x07, 0x2D, 0x74, 0x02, 0x51, 0x5A, 0x3E, 0x09, 0x5F, 0x34, 0x2B,
	0x07, 0x31, 0x1D, 0x32, 0x56, 0x25, 0x1A, 0x09, 0x0E, 0x1B, 0x1D, 0x71,
	0x2A, 0x0B, 0x26, 0x01, 0x18, 0x25, 0x0A, 0x08, 0x59, 0x6D, 0x25, 0x29,
	0x2B, 0x1D, 0x00, 0x25, 0x0C, 0x1F, 0x1D, 0x0F, 0x20, 0x27, 0x02, 0x1A,
	0x2C, 0x3B, 0x12, 0x19, 0x1D, 0x2C, 0x5C, 0x54, 0x26, 0x3A, 0x2A, 0x1B,
	0x52, 0x3E, 0x5B, 0x7B, 0x14, 0x35, 0x20, 0x0E, 0x13, 0x0B, 0x57, 0x58,
	0x44, 0x33, 0x25, 0x18, 0x2A, 0x53, 0x24, 0x26, 0x17, 0x24, 0x5C, 0x69,
	0x34, 0x05, 0x5F, 0x2D, 0x1A, 0x3D, 0x2C, 0x29, 0x32, 0x33, 0x04, 0x0F,
	0x1A, 0x1E, 0x08, 0x25, 0x06, 0x03, 0x0C, 0x36, 0x38, 0x1B, 0x5F, 0x0D,
	0x14, 0x2D, 0x16, 0x59, 0x06, 0x11, 0x08, 0x16, 0x17, 0x07, 0x2D, 0x3E,
	0x03, 0x5B, 0x23, 0x09, 0x3D, 0x2E, 0x27, 0x3F, 0x2A, 0x35, 0x2B, 0x1A,
	0x00, 0x12, 0x5F, 0x51, 0x22, 0x07, 0x04, 0x36, 0x08, 0x05, 0x0E, 0x7B,
	0x54, 0x07, 0x2A, 0x05, 0x2A, 0x5A, 0x28, 0x1C, 0x11, 0x75, 0x54, 0x02,
	0x2B, 0x0A, 0x15, 0x15, 0x02, 0x2D, 0x2E, 0x0D, 0x15, 0x15, 0x28, 0x09,
	0x0F, 0x3B, 0x2B, 0x2D, 0x40, 0x0C, 0x15, 0x0A, 0x25, 0x29, 0x21, 0x19,
	0x23, 0x2C, 0x38, 0x21, 0x3E, 0x58, 0x23, 0x13, 0x24, 0x1E, 0x36, 0x0D,
	0x01, 0x0D, 0x5E, 0x0C, 0x1B, 0x11, 0x07, 0x05, 0x06, 0x59, 0x40, 0x12,
	0x1A, 0x33, 0x5D, 0x2A, 0x0C, 0x5E, 0x35, 0x28, 0x33, 0x72, 0x2D, 0x37,
	0x5F, 0x3D, 0x00, 0x2E, 0x2B, 0x21, 0x29, 0x26, 0x1E, 0x0A, 0x36, 0x06,
	0x34, 0x25, 0x57, 0x58, 0x5D, 0x12, 0x0D, 0x06, 0x2B, 0x08, 0x01, 0x07,
	0x20, 0x16, 0x00, 0x2A, 0x19, 0x2B, 0x5B, 0x05, 0x05, 0x19, 0x38, 0x2A,
	0x5A, 0x0D, 0x20, 0x30, 0x0C, 0x3F, 0x28, 0x2A, 0x31, 0x0C, 0x01, 0x77,
	0x59, 0x17, 0x19, 0x3D, 0x26, 0x36, 0x0C, 0x0D, 0x0D, 0x23, 0x3F, 0x55,
	0x18, 0x09, 0x37, 0x21, 0x37, 0x23, 0x23, 0x18, 0x15, 0x51, 0x09, 0x3D,
	0x0E, 0x21, 0x0E, 0x2F, 0x12, 0x34, 0x5D, 0x53, 0x39, 0x3D, 0x13, 0x34,
	0x07, 0x37, 0x52, 0x0D, 0x59, 0x11, 0x05, 0x0E, 0x2D, 0x0B, 0x15, 0x20,
	0x40, 0x23, 0x09, 0x51, 0x0B, 0x5B, 0x72, 0x18, 0x50, 0x0D, 0x3D, 0x20,
	0x1F, 0x38, 0x5C, 0x38, 0x0C, 0x3F, 0x06, 0x07, 0x26, 0x2E, 0x55, 0x38,
	0x06, 0x04, 0x10, 0x1B, 0x32, 0x3E, 0x2F, 0x2D, 0x08, 0x24, 0x3C, 0x2C,
	0x30, 0x3A, 0x09, 0x23, 0x2C, 0x7A, 0x39, 0x12, 0x5D, 0x2C, 0x3A, 0x38,
	0x0B, 0x2A, 0x53, 0x36, 0x05, 0x59, 0x59, 0x3E, 0x08, 0x00, 0x05, 0x2D,
	0x04, 0x1A, 0x09, 0x36, 0x0F, 0x0E, 0x12, 0x2B, 0x24, 0x5D, 0x1D, 0x18,
	0x25, 0x39, 0x37, 0x27, 0x73, 0x27, 0x32, 0x02, 0x3A, 0x06, 0x19, 0x13,
	0x1D, 0x25, 0x38, 0x5D, 0x32, 0x06, 0x52, 0x73, 0x00, 0x2D, 0x08, 0x44,
	0x0B, 0x0F, 0x2B, 0x37, 0x5A, 0x0A, 0x08, 0x30, 0x3C, 0x12, 0x2C, 0x21,
	0x52, 0x01, 0x5E, 0x2A, 0x5F, 0x12, 0x1E, 0x25, 0x2B, 0x34, 0x3B, 0x28,
	0x3F, 0x0E, 0x0D, 0x05, 0x1F, 0x21, 0x0A, 0x07, 0x05, 0x36, 0x32, 0x7A,
	0x08, 0x28, 0x2C, 0x23, 0x6D, 0x3C, 0x00, 0x5C, 0x24, 0x69, 0x26, 0x39,
	0x2B, 0x08, 0x34, 0x1D, 0x38, 0x25, 0x3C, 0x0F, 0x5A, 0x57, 0x26, 0x13,
	0x1B, 0x27, 0x4E, 0x3D, 0x1D, 0x6D, 0x28, 0x17, 0x59, 0x19, 0x18, 0x02,
	0x56, 0x27, 0x1B, 0x71, 0x54, 0x34, 0x01, 0x32, 0x18, 0x2E, 0x53, 0x09,
	0x20, 0x77, 0x06, 0x20, 0x2F, 0x1A, 0x2C, 0x23, 0x0D, 0x57, 0x2A, 0x2A,
	0x02, 0x0C, 0x45, 0x33, 0x3B, 0x5F, 0x24, 0x56, 0x05, 0x2F, 0x25, 0x2A,
	0x0D, 0x07, 0x2B, 0x06, 0x12, 0x5F, 0x1E, 0x0D, 0x23, 0x23, 0x58, 0x2E,
	0x69, 0x3B, 0x18, 0x2B, 0x5A, 0x25, 0x3C, 0x39, 0x06, 0x06, 0x2A, 0x5F,
	0x54, 0x37, 0x58, 0x28, 0x20, 0x27, 0x17, 0x1D, 0x33, 0x35, 0x50, 0x0B,
	0x33, 0x74, 0x2E, 0x39, 0x16, 0x44, 0x77, 0x2D, 0x28, 0x5A, 0x3E, 0x20,
	0x0F, 0x4A, 0x25, 0x21, 0x7A, 0x28, 0x53, 0x3B, 0x2D, 0x04, 0x38, 0x56,
	0x09, 0x03, 0x75, 0x36, 0x18, 0x0D, 0x2A, 0x69, 0x5F, 0x57, 0x2D, 0x31,
	0x26, 0x34, 0x2F, 0x07, 0x04, 0x15, 0x09, 0x17, 0x5A, 0x21, 0x0A, 0x25,
	0x12, 0x3E, 0x0E, 0x30, 0x01, 0x56, 0x57, 0x2E, 0x20, 0x21, 0x14, 0x0D,
	0x2A, 0x2D, 0x5F, 0x13, 0x09, 0x19, 0x0D, 0x3E, 0x4A, 0x0C, 0x12, 0x08,
	0x3C, 0x2F, 0x0D, 0x5A, 0x24, 0x3F, 0x24, 0x01, 0x3D, 0x36, 0x1F, 0x27,
	0x3F, 0x02, 0x24, 0x18, 0x16, 0x02, 0x19, 0x69, 0x43, 0x10, 0x39, 0x5F,
	0x06, 0x36, 0x34, 0x14, 0x06, 0x05, 0x5A, 0x0F, 0x00, 0x09, 0x76, 0x25,
	0x50, 0x1C, 0x12, 0x04, 0x55, 0x0D, 0x5E, 0x1B, 0x17, 0x07, 0x12, 0x5B,
	0x3F, 0x38, 0x14, 0x33, 0x34, 0x5E, 0x0C, 0x43, 0x24, 0x14, 0x2D, 0x35,
	0x43, 0x12, 0x04, 0x31, 0x0B, 0x06, 0x17, 0x39, 0x32, 0x32, 0x0A, 0x31,
	0x39, 0x2E, 0x34, 0x5E, 0x12, 0x36, 0x01, 0x14, 0x22, 0x37, 0x1F, 0x53,
	0x74, 0x01, 0x24, 0x1A, 0x5F, 0x2E, 0x55, 0x16, 0x2D, 0x40, 0x16, 0x58,
	0x2C, 0x0C, 0x5B, 0x01, 0x28, 0x30, 0x34, 0x3F, 0x70, 0x54, 0x05, 0x0C,
	0x39, 0x72, 0x03, 0x27, 0x0D, 0x25, 0x07, 0x18, 0x50, 0x0D, 0x5C, 0x24,
	0x54, 0x07, 0x09, 0x23, 0x7A, 0x25, 0x53, 0x23, 0x1A, 0x2A, 0x06, 0x0C,
	0x09, 0x5D, 0x04, 0x24, 0x05, 0x27, 0x58, 0x14, 0x07, 0x04, 0x58, 0x01,
	0x2E, 0x28, 0x57, 0x59, 0x2A, 0x1A, 0x09, 0x20, 0x1F, 0x04, 0x0A, 0x22,
	0x08, 0x2B, 0x1A, 0x24, 0x3A, 0x15, 0x00, 0x40, 0x0C, 0x00, 0x2F, 0x23,
	0x1D, 0x2B, 0x27, 0x51, 0x03, 0x3E, 0x3B, 0x5B, 0x19, 0x24, 0x5D, 0x20,
	0x3B, 0x27, 0x04, 0x3D, 0x23, 0x16, 0x06, 0x22, 0x3D, 0x69, 0x29, 0x08,
	0x00, 0x0A, 0x28, 0x0F, 0x17, 0x34, 0x28, 0x2F, 0x35, 0x4E, 0x05, 0x25,
	0x26, 0x2E, 0x2D, 0x27, 0x29, 0x07, 0x1B, 0x11, 0x14, 0x25, 0x76, 0x20,
	0x31, 0x3E, 0x05, 0x04, 0x26, 0x05, 0x1C, 0x59, 0x2D, 0x28, 0x02, 0x00,
	0x0F, 0x72, 0x01, 0x38, 0x5B, 0x1C, 0x0E, 0x09, 0x2F, 0x2F, 0x27, 0x27,
	0x5B, 0x28, 0x18, 0x0C, 0x06, 0x36, 0x13, 0x0D, 0x59, 0x11, 0x2B, 0x56,
	0x5E, 0x01, 0x70, 0x21, 0x2D, 0x02, 0x3E, 0x0F, 0x34, 0x33, 0x1C, 0x44,
	0x06, 0x00, 0x52, 0x23, 0x0C, 0x01, 0x59, 0x17, 0x22, 0x5F, 0x2F, 0x43,
	0x13, 0x58, 0x2A, 0x26, 0x1A, 0x10, 0x2D, 0x01, 0x12, 0x15, 0x3B, 0x3B,
	0x07, 0x72, 0x58, 0x27, 0x26, 0x3F, 0x06, 0x3D, 0x05, 0x01, 0x3E, 0x6D,
	0x0B, 0x20, 0x06, 0x3F, 0x2A, 0x09, 0x24, 0x0B, 0x5A, 0x21, 0x25, 0x12,
	0x26, 0x5B, 0x2D, 0x2F, 0x12, 0x23, 0x3B, 0x05, 0x00, 0x14, 0x26, 0x02,
	0x28, 0x5C, 0x09, 0x3B, 0x3F, 0x00, 0x08, 0x4E, 0x3C, 0x33, 0x04, 0x15,
	0x06, 0x18, 0x18, 0x37, 0x5C, 0x08, 0x03, 0x1E, 0x11, 0x5C, 0x33, 0x56,
	0x40, 0x2D, 0x3F, 0x20, 0x37, 0x3B, 0x2D, 0x1A, 0x39, 0x1E, 0x01, 0x30,
	0x15, 0x13, 0x16, 0x05, 0x01, 0x39, 0x39, 0x1A, 0x04, 0x20, 0x1A, 0x35,
	0x57, 0x2A, 0x30, 0x54, 0x15, 0x1E, 0x58, 0x2D, 0x0E, 0x37, 0x20, 0x1E,
	0x0F, 0x19, 0x2C, 0x3C, 0x22, 0x31, 0x34, 0x55, 0x24, 0x07, 0x77, 0x0F,
	0x57, 0x16, 0x58, 0x20, 0x27, 0x51, 0x1B, 0x3E, 0x16, 0x0A, 0x2E, 0x45,
	0x5A, 0x26, 0x21, 0x59, 0x3E, 0x0D, 0x73, 0x35, 0x51, 0x27, 0x5A, 0x0D,
	0x1F, 0x0A, 0x16, 0x32, 0x09, 0x20, 0x0B, 0x08, 0x32, 0x77, 0x3D, 0x55,
	0x2C, 0x1A, 0x2D, 0x2B, 0x20, 0x1B, 0x39, 0x20, 0x0D, 0x2B, 0x2A, 0x00,
	0x1B, 0x43, 0x29, 0x00, 0x07, 0x37, 0x1C, 0x53, 0x16, 0x59, 0x3A, 0x1D,
	0x08, 0x0A, 0x58, 0x74, 0x3A, 0x20, 0x3C, 0x0E, 0x0B, 0x21, 0x14, 0x28,
	0x5A, 0x72, 0x23, 0x15, 0x00, 0x5B, 0x2B, 0x2D, 0x18, 0x36, 0x5A, 0x11,
	0x2D, 0x0A, 0x5B, 0x12, 0x08, 0x5E, 0x50, 0x28, 0x1A, 0x25, 0x1A, 0x2E,
	0x2C, 0x5F, 0x29, 0x09, 0x57, 0x2B, 0x3B, 0x09, 0x0D, 0x51, 0x3E, 0x04,
	0x04, 0x1C, 0x23, 0x29, 0x13, 0x2C, 0x19, 0x4A, 0x24, 0x0D, 0x77, 0x14,
	0x52, 0x0C, 0x0F, 0x10, 0x43, 0x0D, 0x26, 0x53, 0x20, 0x36, 0x33, 0x41,
	0x58, 0x12, 0x1F, 0x56, 0x56, 0x32, 0x7B, 0x5C, 0x14, 0x03, 0x1A, 0x1A,
	0x16, 0x4E, 0x5A, 0x59, 0x3B, 0x06, 0x59, 0x25, 0x07, 0x0C, 0x3F, 0x03,
	0x18, 0x00, 0x15, 0x47, 0x12, 0x38, 0x58, 0x35, 0x22, 0x29, 0x2F, 0x26,
	0x7A, 0x5A, 0x25, 0x05, 0x22, 0x07, 0x06, 0x35, 0x3B, 0x26, 0x34, 0x36,
	0x2E, 0x5C, 0x01, 0x33, 0x55, 0x23, 0x2F, 0x20, 0x03, 0x20, 0x0A, 0x3C,
	0x28, 0x0E, 0x3E, 0x27, 0x03, 0x32, 0x76, 0x25, 0x50, 0x2D, 0x20, 0x76,
	0x0A, 0x10, 0x22, 0x0C, 0x20, 0x3D, 0x1B, 0x1C, 0x0E, 0x30, 0x25, 0x03,
	0x0F, 0x2E, 0x23, 0x18, 0x57, 0x3E, 0x01, 0x76, 0x02, 0x2E, 0x34, 0x02,
	0x34, 0x2E, 0x56, 0x0F, 0x18, 0x6D, 0x5B, 0x28, 0x3E, 0x29, 0x69, 0x2B,
	0x17, 0x03, 0x02, 0x1A, 0x0A, 0x51, 0x1D, 0x2A, 0x12, 0x1A, 0x2C, 0x41,
	0x2A, 0x34, 0x2D, 0x0E, 0x06, 0x27, 0x71, 0x5B, 0x05, 0x37, 0x21, 0x13,
	0x06, 0x33, 0x5D, 0x22, 0x0B, 0x1B, 0x3B, 0x2D, 0x5D, 0x70, 0x14, 0x50,
	0x18, 0x5E, 0x0F, 0x3B, 0x39, 0x38, 0x20, 0x2F, 0x5B, 0x07, 0x1A, 0x0F,
	0x34, 0x3F, 0x39, 0x19, 0x2C, 0x07, 0x5F, 0x4A, 0x5B, 0x27, 0x7A, 0x03,
	0x10, 0x1E, 0x03, 0x05, 0x20, 0x20, 0x37, 0x26, 0x2F, 0x03, 0x14, 0x25,
	0x59, 0x15, 0x5C, 0x4A, 0x37, 0x0C, 0x13, 0x00, 0x05, 0x23, 0x19, 0x14,
	0x54, 0x36, 0x0A, 0x2A, 0x13, 0x28, 0x1B, 0x5C, 0x23, 0x0A, 0x25, 0x0A,
	0x09, 0x58, 0x71, 0x34, 0x07, 0x59, 0x23, 0x2F, 0x09, 0x23, 0x1B, 0x3E,
	0x2A, 0x27, 0x57, 0x57, 0x40, 0x16, 0x2D, 0x16, 0x58, 0x1C, 0x6D, 0x21,
	0x2E, 0x56, 0x29, 0x12, 0x04, 0x3B, 0x08, 0x18, 0x18, 0x06, 0x22, 0x21,
	0x09, 0x35, 0x34, 0x0C, 0x37, 0x20, 0x34, 0x0E, 0x2A, 0x56, 0x00, 0x16,
	0x2A, 0x08, 0x26, 0x12, 0x0B, 0x55, 0x59, 0x5E, 0x3E, 0x03, 0x38, 0x10,
	0x5E, 0x28, 0x20, 0x26, 0x2E, 0x41, 0x03, 0x12, 0x04, 0x14, 0x5F, 0x2A,
	0x74, 0x47, 0x4A, 0x3D, 0x2E, 0x0E, 0x28, 0x2D, 0x24, 0x40, 0x3A, 0x2D,
	0x35, 0x14, 0x31, 0x04, 0x29, 0x24, 0x41, 0x3E, 0x33, 0x22, 0x17, 0x22,
	0x59, 0x00, 0x39, 0x19, 0x16, 0x33, 0x2A, 0x3A, 0x0E, 0x21, 0x12, 0x71,
	0x35, 0x37, 0x19, 0x40, 0x0B, 0x5F, 0x58, 0x24, 0x27, 0x2D, 0x19, 0x02,
	0x3D, 0x25, 0x77, 0x27, 0x2C, 0x08, 0x05, 0x23, 0x25, 0x3B, 0x06, 0x13,
	0x2B, 0x3C, 0x4E, 0x08, 0x03, 0x12, 0x24, 0x4E, 0x34, 0x09, 0x1B, 0x29,
	0x2D, 0x21, 0x18, 0x33, 0x5C, 0x03, 0x27, 0x24, 0x7A, 0x2E, 0x4A, 0x1E,
	0x3B, 0x0A, 0x20, 0x4A, 0x2C, 0x02, 0x12, 0x00, 0x18, 0x38, 0x03, 0x01,
	0x3F, 0x0A, 0x08, 0x00, 0x0A, 0x5B, 0x12, 0x21, 0x00, 0x20, 0x47, 0x12,
	0x21, 0x29, 0x72, 0x2B, 0x54, 0x3A, 0x29, 0x09, 0x54, 0x10, 0x00, 0x2A,
	0x35, 0x5A, 0x35, 0x1B, 0x5A, 0x25, 0x3D, 0x13, 0x3C, 0x2D, 0x21, 0x2A,
	0x22, 0x2F, 0x09, 0x2C, 0x25, 0x12, 0x0D, 0x5A, 0x05, 0x24, 0x4E, 0x58,
	0x01, 0x20, 0x35, 0x25, 0x3A, 0x19, 0x75, 0x02, 0x1B, 0x59, 0x19, 0x11,
	0x5B, 0x3B, 0x09, 0x52, 0x34, 0x1F, 0x25, 0x27, 0x02, 0x69, 0x26, 0x24,
	0x1A, 0x2F, 0x2D, 0x54, 0x0B, 0x45, 0x28, 0x32, 0x26, 0x07, 0x05, 0x00,
	0x21, 0x2F, 0x57, 0x5F, 0x44, 0x04, 0x3C, 0x08, 0x06, 0x32, 0x7B, 0x47,
	0x06, 0x59, 0x11, 0x35, 0x1A, 0x59, 0x3F, 0x06, 0x38, 0x08, 0x52, 0x01,
	0x18, 0x2B, 0x34, 0x54, 0x29, 0x5C, 0x3B, 0x5C, 0x11, 0x3C, 0x31, 0x72,
	0x1F, 0x24, 0x1B, 0x44, 0x18, 0x0B, 0x02, 0x37, 0x11, 0x25, 0x07, 0x12,
	0x5A, 0x5C, 0x10, 0x58, 0x39, 0x5B, 0x1E, 0x30, 0x28, 0x2B, 0x04, 0x5B,
	0x0C, 0x02, 0x03, 0x5B, 0x21, 0x34, 0x3D, 0x54, 0x28, 0x0C, 0x2D, 0x28,
	0x09, 0x58, 0x0C, 0x05, 0x3C, 0x36, 0x17, 0x39, 0x38, 0x1E, 0x24, 0x22,
	0x06, 0x06, 0x29, 0x22, 0x2C, 0x3C, 0x7B, 0x3E, 0x25, 0x27, 0x3F, 0x18,
	0x2D, 0x11, 0x2C, 0x19, 0x77, 0x27, 0x1B, 0x2D, 0x24, 0x25, 0x35, 0x39,
	0x21, 0x0A, 0x35, 0x14, 0x54, 0x59, 0x02, 0x6D, 0x36, 0x09, 0x1F, 0x11,
	0x38, 0x27, 0x20, 0x07, 0x03, 0x3A, 0x24, 0x1B, 0x25, 0x2E, 0x0E, 0x2A,
	0x27, 0x16, 0x0E, 0x7B, 0x02, 0x55, 0x3A, 0x1F, 0x0F, 0x04, 0x50, 0x22,
	0x29, 0x24, 0x58, 0x0F, 0x45, 0x39, 0x07, 0x1D, 0x07, 0x03, 0x2E, 0x15,
	0x2D, 0x00, 0x21, 0x38, 0x12, 0x03, 0x51, 0x2F, 0x04, 0x73, 0x54, 0x31,
	0x2A, 0x32, 0x1B, 0x24, 0x2E, 0x0B, 0x1F, 0x0D, 0x29, 0x11, 0x0A, 0x3F,
	0x34, 0x15, 0x3B, 0x5D, 0x12, 0x2C, 0x5F, 0x16, 0x37, 0x22, 0x75, 0x54,
	0x14, 0x04, 0x59, 0x72, 0x59, 0x08, 0x02, 0x5D, 0x04, 0x25, 0x2D, 0x27,
	0x44, 0x73, 0x0D, 0x19, 0x1F, 0x53, 0x38, 0x15, 0x13, 0x09, 0x2D, 0x27,
	0x0B, 0x0B, 0x14, 0x1D, 0x27, 0x19, 0x4E, 0x3F, 0x20, 0x0F, 0x43, 0x56,
	0x01, 0x23, 0x0C, 0x36, 0x14, 0x0A, 0x0A, 0x0D, 0x1F, 0x33, 0x05, 0x5F,
	0x3B, 0x55, 0x59, 0x34, 0x53, 0x74, 0x18, 0x10, 0x34, 0x53, 0x20, 0x21,
	0x38, 0x3C, 0x11, 0x7B, 0x2D, 0x02, 0x0F, 0x20, 0x71, 0x1A, 0x0E, 0x25,
	0x11, 0x3B, 0x1D, 0x34, 0x16, 0x1E, 0x36, 0x18, 0x06, 0x18, 0x1D, 0x23,
	0x21, 0x2D, 0x45, 0x33, 0x77, 0x2E, 0x3B, 0x59, 0x13, 0x29, 0x02, 0x02,
	0x1D, 0x39, 0x2B, 0x03, 0x08, 0x0D, 0x12, 0x3B, 0x16, 0x0A, 0x3D, 0x06,
	0x76, 0x23, 0x11, 0x3E, 0x3C, 0x2B, 0x58, 0x35, 0x03, 0x1C, 0x7A, 0x14,
	0x58, 0x04, 0x5C, 0x75, 0x27, 0x54, 0x19, 0x11, 0x21, 0x1D, 0x12, 0x57,
	0x0C, 0x37, 0x08, 0x10, 0x04, 0x39, 0x32, 0x5A, 0x2A, 0x07, 0x09, 0x2A,
	0x21, 0x4A, 0x37, 0x0C, 0x2F, 0x18, 0x02, 0x20, 0x0A, 0x27, 0x2B, 0x11,
	0x1C, 0x53, 0x09, 0x5C, 0x0E, 0x21, 0x2E, 0x69, 0x2D, 0x04, 0x2B, 0x18,
	0x0A, 0x0F, 0x54, 0x1B, 0x27, 0x7B, 0x24, 0x27, 0x56, 0x28, 0x6D, 0x5D,
	0x29, 0x37, 0x07, 0x25, 0x23, 0x05, 0x45, 0x39, 0x01, 0x20, 0x03, 0x56,
	0x13, 0x0B, 0x06, 0x06, 0x29, 0x3F, 0x32, 0x29, 0x56, 0x29, 0x0F, 0x25,
	0x5C, 0x26, 0x5A, 0x2D, 0x15, 0x2E, 0x05, 0x3E, 0x29, 0x0C, 0x03, 0x0D,
	0x2A, 0x33, 0x10, 0x09, 0x55, 0x41, 0x3E, 0x34, 0x35, 0x59, 0x5B, 0x19,
	0x26, 0x24, 0x38, 0x45, 0x3B, 0x76, 0x58, 0x2E, 0x20, 0x29, 0x30, 0x2D,
	0x16, 0x5C, 0x25, 0x3A, 0x08, 0x22, 0x2D, 0x5F, 0x2A, 0x1A, 0x31, 0x0F,
	0x59, 0x12, 0x1E, 0x1B, 0x07, 0x26, 0x69, 0x02, 0x20, 0x18, 0x08, 0x13,
	0x3C, 0x03, 0x2F, 0x25, 0x2D, 0x03, 0x55, 0x1F, 0x3A, 0x23, 0x21, 0x23,
	0x1E, 0x5D, 0x6D, 0x43, 0x0D, 0x29, 0x00, 0x07, 0x3F, 0x20, 0x0D, 0x0D,
	0x05, 0x36, 0x09, 0x2D, 0x18, 0x0D, 0x1D, 0x4E, 0x3C, 0x2A, 0x16, 0x34,
	0x16, 0x59, 0x03, 0x72, 0x2D, 0x03, 0x3A, 0x04, 0x2B, 0x3D, 0x56, 0x29,
	0x53, 0x1A, 0x06, 0x50, 0x58, 0x0D, 0x7A, 0x3B, 0x20, 0x18, 0x28, 0x03,
	0x02, 0x02, 0x59, 0x05, 0x29, 0x35, 0x54, 0x3D, 0x3F, 0x71, 0x15, 0x23,
	0x14, 0x22, 0x0F, 0x35, 0x56, 0x29, 0x31, 0x09, 0x21, 0x00, 0x5C, 0x5F,
	0x2F, 0x3B, 0x04, 0x1D, 0x31, 0x2B, 0x19, 0x59, 0x17, 0x53, 0x77, 0x2A,
	0x0A, 0x00, 0x0D, 0x25, 0x06, 0x2B, 0x5F, 0x5F, 0x24, 0x3A, 0x2C, 0x0B,
	0x07, 0x2F, 0x3A, 0x12, 0x5E, 0x02, 0x75, 0x1A, 0x23, 0x5E, 0x0C, 0x34,
	0x18, 0x29, 0x58, 0x0D, 0x3B, 0x20, 0x29, 0x5A, 0x38, 0x18, 0x1A, 0x32,
	0x2C, 0x39, 0x2A, 0x19, 0x22, 0x01, 0x2E, 0x27, 0x20, 0x4A, 0x38, 0x2A,
	0x23, 0x0B, 0x0C, 0x14, 0x01, 0x7A, 0x5A, 0x14, 0x20, 0x04, 0x2B, 0x2A,
	0x28, 0x3A, 0x1F, 0x0A, 0x2D, 0x0F, 0x2D, 0x53, 0x03, 0x3A, 0x0D, 0x06,
	0x58, 0x72, 0x5B, 0x06, 0x25, 0x27, 0x25, 0x5F, 0x51, 0x25, 0x31, 0x30,
	0x2B, 0x04, 0x09, 0x3B, 0x31, 0x3D, 0x07, 0x58, 0x2F, 0x04, 0x3B, 0x32,
	0x37, 0x1E, 0x3B, 0x5E, 0x22, 0x2F, 0x28, 0x25, 0x06, 0x25, 0x0D, 0x23,
	0x37, 0x58, 0x23, 0x0A, 0x3F, 0x1A, 0x0A, 0x59, 0x38, 0x2E, 0x25, 0x36,
	0x36, 0x5E, 0x3A, 0x17, 0x36, 0x28, 0x08, 0x31, 0x73, 0x36, 0x09, 0x26,
	0x3A, 0x18, 0x2A, 0x29, 0x08, 0x08, 0x09, 0x01, 0x20, 0x2B, 0x2E, 0x0E,
	0x24, 0x19, 0x59, 0x23, 0x15, 0x5C, 0x0C, 0x3E, 0x59, 0x08, 0x3E, 0x2B,
	0x1B, 0x08, 0x01, 0x3D, 0x06, 0x39, 0x59, 0x0B, 0x1E, 0x12, 0x23, 0x5D,
	0x15, 0x24, 0x50, 0x16, 0x3A, 0x0B, 0x22, 0x2F, 0x3A, 0x0C, 0x0B, 0x5A,
	0x0F, 0x5B, 0x3A, 0x0E, 0x3B, 0x11, 0x5A, 0x00, 0x05, 0x5B, 0x4E, 0x45,
	0x29, 0x0D, 0x01, 0x2D, 0x2F, 0x1B, 0x0D, 0x02, 0x55, 0x1F, 0x21, 0x32,
	0x04, 0x52, 0x19, 0x1F, 0x74, 0x14, 0x19, 0x18, 0x59, 0x12, 0x2D, 0x2E,
	0x2B, 0x0D, 0x1A, 0x1F, 0x17, 0x5C, 0x38, 0x0C, 0x47, 0x3B, 0x24, 0x02,
	0x09, 0x1A, 0x0A, 0x07, 0x5C, 0x2C, 0x14, 0x0E, 0x26, 0x23, 0x7A, 0x07,
	0x12, 0x17, 0x22, 0x2D, 0x14, 0x12, 0x0F, 0x13, 0x70, 0x2E, 0x37, 0x2A,
	0x27, 0x17, 0x58, 0x0B, 0x37, 0x26, 0x0A, 0x5B, 0x07, 0x39, 0x13, 0x3B,
	0x0E, 0x03, 0x2F, 0x39, 0x77, 0x47, 0x2C, 0x1F, 0x3F, 0x75, 0x3F, 0x37,
	0x00, 0x2C, 0x0E, 0x5E, 0x1B, 0x0B, 0x1E, 0x72, 0x2D, 0x50, 0x1B, 0x29,
	0x17, 0x3B, 0x39, 0x3D, 0x19, 0x3A, 0x0B, 0x29, 0x21, 0x59, 0x05, 0x04,
	0x1B, 0x38, 0x22, 0x2A, 0x09, 0x2B, 0x5A, 0x02, 0x0C, 0x47, 0x35, 0x09,
	0x11, 0x6D, 0x3B, 0x02, 0x36, 0x05, 0x07, 0x19, 0x24, 0x1A, 0x13, 0x1A,
	0x08, 0x34, 0x28, 0x3B, 0x2C, 0x3B, 0x03, 0x58, 0x23, 0x12, 0x0B, 0x02,
	0x19, 0x33, 0x0C, 0x34, 0x36, 0x07, 0x27, 0x2A, 0x28, 0x2F, 0x5B, 0x39,
	0x20, 0x00, 0x2E, 0x3D, 0x5B, 0x29, 0x38, 0x17, 0x3D, 0x13, 0x13, 0x16,
	0x03, 0x25, 0x00, 0x32, 0x02, 0x08, 0x34, 0x5E, 0x30, 0x35, 0x0F, 0x01,
	0x0E, 0x17, 0x03, 0x26, 0x2F, 0x22, 0x36, 0x55, 0x00, 0x5E, 0x33, 0x1A,
	0x5B, 0x11, 0x03, 0x38, 0x26, 0x5E, 0x55, 0x20, 0x5E, 0x25, 0x0A, 0x56,
	0x06, 0x08, 0x24, 0x3C, 0x56, 0x2D, 0x33, 0x2F, 0x09, 0x52, 0x3E, 0x32,
	0x20, 0x24, 0x0B, 0x0A, 0x02, 0x0C, 0x25, 0x2D, 0x22, 0x5C, 0x07, 0x5A,
	0x08, 0x23, 0x08, 0x26, 0x2B, 0x59, 0x3E, 0x59, 0x04, 0x2F, 0x06, 0x5A,
	0x38, 0x2F, 0x54, 0x59, 0x27, 0x23, 0x10, 0x35, 0x2A, 0x5D, 0x1A, 0x27,
	0x38, 0x34, 0x03, 0x06, 0x72, 0x1C, 0x22, 0x5C, 0x27, 0x24, 0x04, 0x35,
	0x57, 0x27, 0x75, 0x0E, 0x00, 0x04, 0x04, 0x71, 0x35, 0x17, 0x23, 0x40,
	0x01, 0x55, 0x11, 0x22, 0x0C, 0x76, 0x5F, 0x19, 0x21, 0x3D, 0x37, 0x00,
	0x57, 0x5C, 0x44, 0x0F, 0x21, 0x33, 0x37, 0x1F, 0x2C, 0x24, 0x07, 0x04,
	0x2F, 0x2A, 0x5D, 0x0F, 0x1D, 0x5E, 0x35, 0x2B, 0x34, 0x3B, 0x03, 0x21,
	0x25, 0x0C, 0x41, 0x1F, 0x18, 0x47, 0x19, 0x2F, 0x1C, 0x10, 0x5F, 0x2C,
	0x23, 0x00, 0x31, 0x02, 0x18, 0x19, 0x12, 0x07, 0x47, 0x28, 0x1D, 0x22,
	0x23, 0x09, 0x25, 0x5D, 0x26, 0x15, 0x0E, 0x3B, 0x16, 0x23, 0x1A, 0x14,
	0x3B, 0x1A, 0x07, 0x34, 0x01, 0x0D, 0x03, 0x59, 0x2D, 0x3A, 0x2E, 0x14,
	0x5C, 0x01, 0x08, 0x0C, 0x02, 0x04, 0x15, 0x0F, 0x4E, 0x5F, 0x3C, 0x0F,
	0x5D, 0x3B, 0x45, 0x02, 0x24, 0x55, 0x4E, 0x16, 0x24, 0x0C, 0x1E, 0x4E,
	0x00, 0x5A, 0x07, 0x1B, 0x51, 0x5B, 0x1E, 0x24, 0x07, 0x30, 0x5C, 0x59,
	0x00, 0x54, 0x0F, 0x3E, 0x40, 0x72, 0x27, 0x28, 0x19, 0x19, 0x0C, 0x02,
	0x55, 0x1D, 0x24, 0x2F, 0x27, 0x59, 0x1A, 0x2C, 0x0D, 0x08, 0x24, 0x0A,
	0x40, 0x16, 0x00, 0x06, 0x3D, 0x58, 0x05, 0x0D, 0x14, 0x3E, 0x11, 0x0D,
	0x2A, 0x59, 0x18, 0x40, 0x16, 0x20, 0x4E, 0x1C, 0x39, 0x20, 0x5D, 0x0A,
	0x2F, 0x3D, 0x71, 0x1A, 0x07, 0x14, 0x28, 0x28, 0x5C, 0x37, 0x59, 0x2F,
	0x3B, 0x15, 0x08, 0x22, 0x2F, 0x06, 0x22, 0x27, 0x08, 0x5D, 0x0C, 0x09,
	0x31, 0x26, 0x2E, 0x17, 0x5D, 0x2B, 0x27, 0x5E, 0x0D, 0x0B, 0x0E, 0x2F,
	0x0E, 0x31, 0x1D, 0x29, 0x14, 0x3B, 0x71, 0x09, 0x35, 0x5D, 0x23, 0x0A,
	0x5F, 0x14, 0x09, 0x19, 0x32, 0x09, 0x22, 0x16, 0x5D, 0x18, 0x54, 0x32,
	0x1F, 0x5E, 0x6D, 0x5F, 0x10, 0x0B, 0x31, 0x2F, 0x19, 0x18, 0x07, 0x29,
	0x0A, 0x3A, 0x29, 0x21, 0x20, 0x07, 0x22, 0x17, 0x06, 0x5D, 0x2C, 0x18,
	0x23, 0x1E, 0x5D, 0x16, 0x47, 0x03, 0x02, 0x3A, 0x73, 0x02, 0x37, 0x3D,
	0x27, 0x75, 0x05, 0x07, 0x37, 0x5A, 0x6D, 0x0B, 0x0C, 0x3E, 0x24, 0x32,
	0x02, 0x15, 0x2C, 0x2A, 0x73, 0x3C, 0x26, 0x3E, 0x0A, 0x6D, 0x3B, 0x09,
	0x06, 0x21, 0x06, 0x2E, 0x31, 0x41, 0x00, 0x32, 0x19, 0x17, 0x2A, 0x0D,
	0x09, 0x3B, 0x37, 0x26, 0x1D, 0x11, 0x1A, 0x54, 0x39, 0x5C, 0x14, 0x0A,
	0x0E, 0x26, 0x1C, 0x7B, 0x0B, 0x22, 0x38, 0x5D, 0x7A, 0x3E, 0x2C, 0x45,
	0x31, 0x26, 0x1F, 0x3B, 0x03, 0x39, 0x11, 0x1F, 0x30, 0x3D, 0x0F, 0x0C,
	0x1B, 0x4E, 0x18, 0x5E, 0x27, 0x2A, 0x27, 0x23, 0x0C, 0x70, 0x0E, 0x16,
	0x41, 0x1B, 0x70, 0x05, 0x36, 0x2C, 0x07, 0x76, 0x04, 0x29, 0x02, 0x1C,
	0x05, 0x06, 0x55, 0x20, 0x53, 0x69, 0x0A, 0x13, 0x5B, 0x0A, 0x0A, 0x1C,
	0x06, 0x0C, 0x2E, 0x36, 0x1C, 0x26, 0x07, 0x20, 0x6D, 0x5A, 0x33, 0x01,
	0x3D, 0x25, 0x35, 0x14, 0x21, 0x5B, 0x1A, 0x5D, 0x32, 0x14, 0x5F, 0x0C,
	0x0F, 0x54, 0x5D, 0x19, 0x77, 0x38, 0x54, 0x34, 0x0C, 0x24, 0x5A, 0x0F,
	0x25, 0x22, 0x2B, 0x0F, 0x50, 0x2F, 0x3B, 0x00, 0x0A, 0x32, 0x2B, 0x19,
	0x21, 0x16, 0x04, 0x3B, 0x28, 0x24, 0x3E, 0x15, 0x24, 0x39, 0x1A, 0x2E,
	0x2C, 0x3B, 0x01, 0x2A, 0x28, 0x52, 0x5D, 0x22, 0x36, 0x2D, 0x2E, 0x3E,
	0x11, 0x71, 0x01, 0x2B, 0x1E, 0x03, 0x2A, 0x54, 0x58, 0x04, 0x5C, 0x3A,
	0x14, 0x2A, 0x1D, 0x40, 0x10, 0x36, 0x56, 0x5A, 0x2C, 0x34, 0x21, 0x2C,
	0x2A, 0x32, 0x2D, 0x0E, 0x36, 0x18, 0x28, 0x1A, 0x0A, 0x1B, 0x03, 0x11,
	0x76, 0x2E, 0x02, 0x06, 0x5B, 0x76, 0x01, 0x27, 0x2F, 0x3B, 0x0E, 0x2F,
	0x23, 0x37, 0x23, 0x25, 0x25, 0x37, 0x07, 0x1F, 0x2C, 0x23, 0x0F, 0x3F,
	0x23, 0x38, 0x20, 0x14, 0x0A, 0x5D, 0x2A, 0x08, 0x55, 0x17, 0x31, 0x25,
	0x3F, 0x32, 0x1B, 0x31, 0x21, 0x58, 0x02, 0x18, 0x3A, 0x3B, 0x5B, 0x18,
	0x5F, 0x40, 0x71, 0x36, 0x14, 0x18, 0x33, 0x3A, 0x27, 0x00, 0x03, 0x1B,
	0x20, 0x14, 0x27, 0x3A, 0x0F, 0x28, 0x47, 0x2A, 0x38, 0x40, 0x37, 0x36,
	0x04, 0x07, 0x1C, 0x29, 0x55, 0x53, 0x00, 0x5D, 0x15, 0x5F, 0x33, 0x24,
	0x07, 0x18, 0x1D, 0x38, 0x36, 0x3E, 0x73, 0x04, 0x0B, 0x19, 0x0A, 0x7A,
	0x04, 0x02, 0x59, 0x31, 0x09, 0x5B, 0x22, 0x3C, 0x27, 0x01, 0x59, 0x0C,
	0x28, 0x5A, 0x7B, 0x38, 0x13, 0x0B, 0x24, 0x05, 0x06, 0x34, 0x02, 0x5B,
	0x0A, 0x0B, 0x27, 0x39, 0x3B, 0x2A, 0x04, 0x57, 0x1F, 0x18, 0x2B, 0x43,
	0x32, 0x03, 0x3B, 0x2C, 0x5B, 0x0C, 0x16, 0x1A, 0x74, 0x58, 0x00, 0x28,
	0x5D, 0x09, 0x29, 0x18, 0x59, 0x09, 0x1A, 0x28, 0x02, 0x2D, 0x1F, 0x2D,
	0x38, 0x18, 0x2D, 0x01, 0x2E, 0x0A, 0x3B, 0x01, 0x58, 0x2F, 0x16, 0x35,
	0x0D, 0x3C, 0x30, 0x23, 0x25, 0x58, 0x2A, 0x07, 0x1C, 0x56, 0x3A, 0x38,
	0x3A, 0x1F, 0x57, 0x25, 0x2F, 0x7B, 0x06, 0x4A, 0x01, 0x5C, 0x37, 0x5A,
	0x0C, 0x3D, 0x32, 0x3A, 0x2D, 0x22, 0x0F, 0x03, 0x20, 0x3D, 0x05, 0x58,
	0x3F, 0x23, 0x0A, 0x4E, 0x5C, 0x59, 0x76, 0x3B, 0x53, 0x1D, 0x31, 0x2F,
	0x26, 0x2F, 0x1C, 0x25, 0x17, 0x2E, 0x3B, 0x37, 0x5B, 0x0B, 0x1B, 0x05,
	0x59, 0x05, 0x3B, 0x3C, 0x54, 0x16, 0x3F, 0x16, 0x5A, 0x0A, 0x56, 0x22,
	0x24, 0x38, 0x05, 0x45, 0x3A, 0x2C, 0x18, 0x16, 0x5B, 0x1C, 0x04, 0x08,
	0x30, 0x2F, 0x52, 0x20, 0x58, 0x34, 0x5E, 0x1E, 0x14, 0x5C, 0x15, 0x41,
	0x21, 0x0D, 0x28, 0x17, 0x45, 0x04, 0x11, 0x19, 0x2D, 0x58, 0x2F, 0x75,
	0x3C, 0x3B, 0x3A, 0x53, 0x10, 0x2D, 0x18, 0x3F, 0x0C, 0x69, 0x02, 0x58,
	0x2F, 0x39, 0x38, 0x55, 0x28, 0x04, 0x18, 0x2A, 0x0A, 0x38, 0x1F, 0x0F,
	0x35, 0x26, 0x20, 0x2C, 0x07, 0x16, 0x23, 0x2E, 0x28, 0x5A, 0x3A, 0x05,
	0x0F, 0x27, 0x07, 0x36, 0x34, 0x12, 0x25, 0x44, 0x00, 0x2D, 0x58, 0x38,
	0x40, 0x2A, 0x29, 0x4E, 0x5D, 0x09, 0x00, 0x2D, 0x31, 0x03, 0x0A, 0x14,
	0x2B, 0x59, 0x25, 0x33, 0x3B, 0x0E, 0x2B, 0x2F, 0x44, 0x3A, 0x2A, 0x38,
	0x18, 0x2E, 0x3B, 0x55, 0x23, 0x2F, 0x04, 0x07, 0x1E, 0x2A, 0x04, 0x0E,
	0x08, 0x43, 0x22, 0x41, 0x38, 0x16, 0x14, 0x28, 0x22, 0x27, 0x7A, 0x03,
	0x31, 0x59, 0x5F, 0x21, 0x22, 0x2B, 0x0F, 0x05, 0x34, 0x22, 0x0B, 0x58,
	0x1E, 0x0D, 0x3B, 0x53, 0x2A, 0x3B, 0x38, 0x5E, 0x32, 0x06, 0x5A, 0x0F,
	0x38, 0x2C, 0x1F, 0x04, 0x04, 0x3E, 0x2F, 0x23, 0x44, 0x34, 0x55, 0x26,
	0x14, 0x19, 0x00, 0x1F, 0x04, 0x04, 0x44, 0x2F, 0x28, 0x2C, 0x1A, 0x27,
	0x06, 0x38, 0x10, 0x37, 0x5B, 0x0E, 0x0A, 0x17, 0x0A, 0x58, 0x33, 0x2B,
	0x33, 0x0C, 0x21, 0x17, 0x2F, 0x32, 0x41, 0x3F, 0x08, 0x5D, 0x3B, 0x5A,
	0x04, 0x77, 0x09, 0x33, 0x00, 0x5D, 0x27, 0x29, 0x07, 0x21, 0x29, 0x04,
	0x5D, 0x28, 0x37, 0x13, 0x27, 0x2D, 0x03, 0x2F, 0x44, 0x0D, 0x58, 0x31,
	0x3D, 0x25, 0x08, 0x16, 0x31, 0x19, 0x32, 0x29, 0x0A, 0x30, 0x2F, 0x11,
	0x17, 0x47, 0x52, 0x18, 0x18, 0x6D, 0x3B, 0x4A, 0x1C, 0x32, 0x2E, 0x2D,
	0x17, 0x08, 0x38, 0x6D, 0x21, 0x00, 0x2C, 0x40, 0x74, 0x09, 0x2F, 0x41,
	0x29, 0x06, 0x39, 0x1B, 0x59, 0x3F, 0x72, 0x28, 0x0C, 0x56, 0x01, 0x75,
	0x47, 0x02, 0x36, 0x23, 0x2F, 0x1A, 0x05, 0x14, 0x5C, 0x6D, 0x2A, 0x30,
	0x3D, 0x27, 0x71, 0x1F, 0x30, 0x3C, 0x5B, 0x1A, 0x0F, 0x2B, 0x28, 0x23,
	0x3A, 0x06, 0x06, 0x5B, 0x1F, 0x2E, 0x5F, 0x2D, 0x3E, 0x5C, 0x21, 0x0E,
	0x4A, 0x2F, 0x2A, 0x28, 0x3F, 0x24, 0x5D, 0x27, 0x04, 0x18, 0x2D, 0x3F,
	0x0D, 0x23, 0x08, 0x09, 0x58, 0x23, 0x37, 0x47, 0x23, 0x14, 0x03, 0x69,
	0x04, 0x36, 0x59, 0x33, 0x77, 0x09, 0x39, 0x27, 0x1C, 0x2D, 0x2F, 0x31,
	0x3F, 0x38, 0x12, 0x2D, 0x12, 0x36, 0x09, 0x2A, 0x0F, 0x39, 0x25, 0x5E,
	0x00, 0x04, 0x0A, 0x1D, 0x1D, 0x2A, 0x58, 0x2F, 0x36, 0x22, 0x15, 0x07,
	0x22, 0x26, 0x1B, 0x27, 0x2B, 0x31, 0x26, 0x33, 0x24, 0x1D, 0x35, 0x00,
	0x1F, 0x0A, 0x5C, 0x26, 0x08, 0x5C, 0x13, 0x0A, 0x16, 0x26, 0x5C, 0x01,
	0x09, 0x30, 0x2A, 0x52, 0x0B, 0x03, 0x35, 0x26, 0x5A, 0x1A, 0x05, 0x22,
	0x0D, 0x24, 0x32, 0x2B, 0x29, 0x3C, 0x0E, 0x6D, 0x43, 0x19, 0x1E, 0x11,
	0x34, 0x5E, 0x31, 0x24, 0x39, 0x77, 0x24, 0x28, 0x0F, 0x33, 0x2F, 0x06,
	0x0A, 0x25, 0x27, 0x75, 0x23, 0x53, 0x0D, 0x5A, 0x71, 0x1F, 0x17, 0x3F,
	0x5C, 0x27, 0x22, 0x2E, 0x59, 0x06, 0x15, 0x1B, 0x19, 0x3E, 0x1E, 0x31,
	0x08, 0x55, 0x24, 0x1E, 0x29, 0x2D, 0x30, 0x1D, 0x1A, 0x0A, 0x5E, 0x0E,
	0x00, 0x1D, 0x03, 0x54, 0x52, 0x01, 0x03, 0x0C, 0x26, 0x58, 0x37, 0x52,
	0x16, 0x5E, 0x2C, 0x3F, 0x03, 0x27, 0x02, 0x25, 0x57, 0x40, 0x28, 0x25,
	0x55, 0x0C, 0x58, 0x2D, 0x59, 0x27, 0x0C, 0x2C, 0x18, 0x22, 0x0A, 0x19,
	0x28, 0x2B, 0x00, 0x0F, 0x5D, 0x00, 0x21, 0x29, 0x32, 0x01, 0x3B, 0x14,
	0x5D, 0x32, 0x09, 0x22, 0x11, 0x55, 0x02, 0x25, 0x12, 0x6D, 0x1D, 0x2C,
	0x2B, 0x1E, 0x15, 0x18, 0x34, 0x1C, 0x0F, 0x09, 0x07, 0x2C, 0x39, 0x00,
	0x6D, 0x2A, 0x30, 0x3C, 0x2E, 0x06, 0x2E, 0x51, 0x2B, 0x1E, 0x1B, 0x20,
	0x3B, 0x03, 0x5C, 0x01, 0x55, 0x05, 0x5A, 0x28, 0x0E, 0x18, 0x4A, 0x03,
	0x0C, 0x00, 0x05, 0x12, 0x0D, 0x32, 0x35, 0x39, 0x54, 0x3C, 0x11, 0x32,
	0x03, 0x53, 0x07, 0x5B, 0x0F, 0x0F, 0x00, 0x0A, 0x07, 0x69, 0x14, 0x29,
	0x3D, 0x22, 0x14, 0x5F, 0x52, 0x5A, 0x40, 0x08, 0x03, 0x2D, 0x21, 0x2A,
	0x32, 0x35, 0x06, 0x1C, 0x2D, 0x06, 0x29, 0x36, 0x2A, 0x3D, 0x31, 0x28,
	0x34, 0x58, 0x27, 0x2C, 0x06, 0x2D, 0x1C, 0x3D, 0x03, 0x27, 0x26, 0x5E,
	0x0D, 0x23, 0x05, 0x0F, 0x25, 0x12, 0x0B, 0x14, 0x4E, 0x20, 0x1E, 0x14,
	0x06, 0x53, 0x2B, 0x11, 0x0B, 0x0F, 0x02, 0x26, 0x04, 0x34, 0x0A, 0x00,
	0x34, 0x2E, 0x16, 0x20, 0x36, 0x39, 0x0E, 0x1B, 0x27, 0x07, 0x20, 0x2C,
	0x04, 0x16, 0x2A, 0x1C, 0x1E, 0x71, 0x47, 0x24, 0x27, 0x3F, 0x2F, 0x26,
	0x29, 0x59, 0x20, 0x13, 0x02, 0x27, 0x21, 0x32, 0x04, 0x58, 0x56, 0x5D,
	0x1B, 0x30, 0x06, 0x14, 0x19, 0x26, 0x11, 0x58, 0x56, 0x5D, 0x53, 0x03,
	0x3B, 0x35, 0x58, 0x28, 0x10, 0x01, 0x0F, 0x5B, 0x2E, 0x2E, 0x3E, 0x23,
	0x58, 0x0D, 0x31, 0x06, 0x05, 0x41, 0x11, 0x7B, 0x16, 0x06, 0x0C, 0x5E,
	0x13, 0x47, 0x3B, 0x45, 0x40, 0x06, 0x0A, 0x4A, 0x05, 0x22, 0x77, 0x14,
	0x57, 0x14, 0x02, 0x17, 0x09, 0x04, 0x14, 0x5F, 0x23, 0x23, 0x30, 0x59,
	0x21, 0x0E, 0x1F, 0x4A, 0x2F, 0x0D, 0x73, 0x24, 0x2C, 0x08, 0x5C, 0x2C,
	0x2D, 0x19, 0x3C, 0x29, 0x38, 0x02, 0x53, 0x07, 0x19, 0x04, 0x25, 0x0A,
	0x3C, 0x2D, 0x21, 0x18, 0x0A, 0x25, 0x28, 0x2B, 0x34, 0x07, 0x28, 0x01,
	0x12, 0x55, 0x2C, 0x38, 0x2A, 0x70, 0x35, 0x29, 0x07, 0x3B, 0x38, 0x0E,
	0x0A, 0x09, 0x05, 0x37, 0x1B, 0x20, 0x09, 0x28, 0x01, 0x04, 0x36, 0x1C,
	0x32, 0x03, 0x0A, 0x16, 0x23, 0x06, 0x32, 0x03, 0x14, 0x5F, 0x18, 0x0A,
	0x2D, 0x13, 0x23, 0x1E, 0x21, 0x2D, 0x59, 0x28, 0x53, 0x00, 0x43, 0x4E,
	0x09, 0x23, 0x06, 0x54, 0x55, 0x2F, 0x05, 0x03, 0x54, 0x05, 0x2C, 0x12,
	0x35, 0x21, 0x29, 0x2A, 0x08, 0x24, 0x0A, 0x15, 0x06, 0x44, 0x07, 0x3C,
	0x04, 0x28, 0x01, 0x06, 0x47, 0x18, 0x3C, 0x5B, 0x0A, 0x35, 0x2E, 0x2F,
	0x0C, 0x3B, 0x5D, 0x4A, 0x06, 0x58, 0x2B, 0x07, 0x02, 0x16, 0x20, 0x35,
	0x1C, 0x54, 0x27, 0x3B, 0x11, 0x27, 0x03, 0x21, 0x40, 0x25, 0x2D, 0x37,
	0x09, 0x2F, 0x2E, 0x0F, 0x28, 0x5A, 0x0C, 0x73, 0x3F, 0x50, 0x36, 0x39,
	0x3A, 0x3C, 0x3B, 0x08, 0x0F, 0x03, 0x2F, 0x0C, 0x05, 0x3A, 0x0F, 0x0D,
	0x3B, 0x1F, 0x21, 0x2D, 0x5E, 0x37, 0x05, 0x5B, 0x05, 0x22, 0x32, 0x38,
	0x0D, 0x2C, 0x34, 0x55, 0x21, 0x32, 0x12, 0x21, 0x22, 0x45, 0x0D, 0x30,
	0x5A, 0x39, 0x1D, 0x04, 0x11, 0x0B, 0x4E, 0x3C, 0x08, 0x30, 0x27, 0x0E,
	0x1B, 0x59, 0x25, 0x26, 0x27, 0x3E, 0x25, 0x33, 0x00, 0x1B, 0x3E, 0x00,
	0x35, 0x21, 0x00, 0x17, 0x13, 0x24, 0x18, 0x08, 0x5E, 0x28, 0x0F, 0x0A,
	0x37, 0x1F, 0x5C, 0x24, 0x23, 0x19, 0x3F, 0x31, 0x34, 0x16, 0x25, 0x01,
	0x31, 0x34, 0x1F, 0x56, 0x5E, 0x22, 0x36, 0x1E, 0x05, 0x19, 0x1F, 0x73,
	0x2D, 0x56, 0x5F, 0x31, 0x74, 0x03, 0x0E, 0x5D, 0x02, 0x3B, 0x59, 0x07,
	0x23, 0x02, 0x38, 0x5C, 0x51, 0x08, 0x0F, 0x10, 0x28, 0x4E, 0x3B, 0x3D,
	0x7B, 0x35, 0x39, 0x1E, 0x24, 0x14, 0x18, 0x09, 0x0B, 0x04, 0x72, 0x0A,
	0x28, 0x38, 0x53, 0x69, 0x5B, 0x16, 0x5D, 0x12, 0x07, 0x18, 0x02, 0x06,
	0x3C, 0x77, 0x26, 0x35, 0x2B, 0x26, 0x21, 0x39, 0x17, 0x09, 0x21, 0x24,
	0x21, 0x13, 0x0C, 0x03, 0x08, 0x36, 0x10, 0x16, 0x05, 0x3B, 0x3D, 0x0E,
	0x5E, 0x3B, 0x18, 0x28, 0x15, 0x24, 0x59, 0x13, 0x20, 0x29, 0x0C, 0x12,
	0x75, 0x47, 0x54, 0x58, 0x3B, 0x03, 0x3F, 0x20, 0x3B, 0x58, 0x09, 0x3A,
	0x05, 0x58, 0x3D, 0x69, 0x2D, 0x32, 0x07, 0x33, 0x2A, 0x0D, 0x04, 0x39,
	0x2A, 0x14, 0x21, 0x03, 0x36, 0x04, 0x36, 0x27, 0x57, 0x3B, 0x2F, 0x3A,
	0x3A, 0x39, 0x5F, 0x00, 0x1A, 0x1C, 0x2B, 0x02, 0x2D, 0x7A, 0x14, 0x13,
	0x17, 0x24, 0x2C, 0x58, 0x04, 0x39, 0x3D, 0x32, 0x18, 0x59, 0x26, 0x2D,
	0x2C, 0x2D, 0x4A, 0x5A, 0x39, 0x13, 0x23, 0x55, 0x04, 0x3A, 0x75, 0x01,
	0x35, 0x1C, 0x53, 0x0D, 0x1B, 0x57, 0x0C, 0x13, 0x75, 0x03, 0x13, 0x1A,
	0x0F, 0x2F, 0x47, 0x07, 0x1D, 0x5F, 0x00, 0x36, 0x39, 0x0B, 0x40, 0x14,
	0x09, 0x0E, 0x36, 0x2E, 0x07, 0x43, 0x39, 0x07, 0x0C, 0x0A, 0x20, 0x03,
	0x2F, 0x27, 0x6D, 0x03, 0x05, 0x0C, 0x2C, 0x28, 0x5E, 0x52, 0x59, 0x29,
	0x6D, 0x38, 0x54, 0x39, 0x0F, 0x38, 0x34, 0x11, 0x3C, 0x27, 0x2F, 0x09,
	0x4E, 0x28, 0x2D, 0x15, 0x1A, 0x26, 0x2A, 0x23, 0x2F, 0x16, 0x2F, 0x1F,
	0x22, 0x1B, 0x26, 0x09, 0x08, 0x0D, 0x04, 0x03, 0x27, 0x03, 0x0F, 0x2B,
	0x1D, 0x33, 0x0A, 0x0E, 0x0E, 0x07, 0x31, 0x5F, 0x5D, 0x3A, 0x3A, 0x4E,
	0x5A, 0x01, 0x2D, 0x02, 0x39, 0x45, 0x01, 0x70, 0x23, 0x30, 0x0F, 0x39,
	0x2E, 0x08, 0x07, 0x39, 0x11, 0x29, 0x3B, 0x1B, 0x3E, 0x52, 0x77, 0x2A,
	0x2C, 0x5D, 0x3A, 0x0E, 0x19, 0x19, 0x01, 0x31, 0x73, 0x5F, 0x00, 0x02,
	0x20, 0x69, 0x55, 0x50, 0x39, 0x2F, 0x72, 0x08, 0x19, 0x1E, 0x44, 0x0E,
	0x28, 0x39, 0x5F, 0x52, 0x29, 0x18, 0x04, 0x5A, 0x5F, 0x73, 0x03, 0x04,
	0x27, 0x0E, 0x2A, 0x1D, 0x39, 0x27, 0x59, 0x3A, 0x58, 0x18, 0x28, 0x3F,
	0x73, 0x3E, 0x12, 0x3B, 0x24, 0x06, 0x59, 0x26, 0x2F, 0x5D, 0x21, 0x5D,
	0x02, 0x1F, 0x53, 0x36, 0x54, 0x20, 0x5C, 0x1D, 0x23, 0x09, 0x0D, 0x59,
	0x21, 0x05, 0x26, 0x57, 0x3B, 0x59, 0x01, 0x09, 0x18, 0x2B, 0x52, 0x04,
	0x0A, 0x10, 0x07, 0x26, 0x0E, 0x39, 0x15, 0x05, 0x5A, 0x77, 0x5C, 0x0A,
	0x23, 0x38, 0x31, 0x1B, 0x08, 0x5D, 0x5B, 0x69, 0x3F, 0x2A, 0x1B, 0x1E,
	0x7A, 0x0E, 0x26, 0x3F, 0x5D, 0x1B, 0x03, 0x27, 0x24, 0x2A, 0x73, 0x5B,
	0x2F, 0x21, 0x1F, 0x13, 0x3F, 0x3B, 0x3D, 0x3C, 0x29, 0x04, 0x20, 0x08,
	0x29, 0x05, 0x54, 0x10, 0x57, 0x12, 0x07, 0x09, 0x20, 0x2F, 0x44, 0x1A,
	0x29, 0x24, 0x23, 0x2F, 0x0E, 0x5F, 0x4A, 0x0A, 0x5E, 0x6D, 0x5B, 0x14,
	0x08, 0x2D, 0x34, 0x26, 0x16, 0x3B, 0x38, 0x0F, 0x1A, 0x2B, 0x2A, 0x33,
	0x09, 0x54, 0x38, 0x0A, 0x09, 0x77, 0x26, 0x04, 0x0F, 0x5A, 0x18, 0x21,
	0x2A, 0x57, 0x53, 0x29, 0x3E, 0x0F, 0x0D, 0x59, 0x05, 0x2E, 0x02, 0x5D,
	0x01, 0x0F, 0x38, 0x03, 0x3F, 0x26, 0x31, 0x2A, 0x25, 0x16, 0x5E, 0x76,
	0x2F, 0x4A, 0x56, 0x1D, 0x18, 0x54, 0x54, 0x41, 0x05, 0x20, 0x5B, 0x2B,
	0x1D, 0x29, 0x16, 0x2B, 0x0A, 0x0A, 0x5B, 0x31, 0x09, 0x33, 0x57, 0x22,
	0x05, 0x15, 0x16, 0x1E, 0x24, 0x11, 0x03, 0x0D, 0x5B, 0x1F, 0x70, 0x5F,
	0x06, 0x2F, 0x44, 0x24, 0x01, 0x1B, 0x05, 0x5D, 0x15, 0x36, 0x2B, 0x5D,
	0x03, 0x71, 0x5B, 0x23, 0x25, 0x44, 0x08, 0x20, 0x11, 0x1F, 0x3E, 0x0C,
	0x1C, 0x08, 0x56, 0x26, 0x27, 0x23, 0x08, 0x45, 0x0E, 0x31, 0x05, 0x18,
	0x06, 0x05, 0x75, 0x2E, 0x20, 0x26, 0x5B, 0x30, 0x05, 0x2E, 0x14, 0x13,
	0x01, 0x3D, 0x23, 0x39, 0x3F, 0x09, 0x23, 0x2D, 0x16, 0x1A, 0x70, 0x04,
	0x2D, 0x0D, 0x0C, 0x0E, 0x22, 0x0A, 0x0C, 0x20, 0x20, 0x0F, 0x36, 0x3E,
	0x28, 0x11, 0x2D, 0x2A, 0x5F, 0x12, 0x09, 0x2A, 0x11, 0x00, 0x5D, 0x03,
	0x27, 0x29, 0x14, 0x05, 0x23, 0x55, 0x06, 0x22, 0x1C, 0x21, 0x21, 0x56,
	0x3F, 0x40, 0x26, 0x1D, 0x51, 0x5E, 0x5A, 0x08, 0x00, 0x2F, 0x1B, 0x28,
	0x21, 0x47, 0x0D, 0x59, 0x38, 0x2F, 0x18, 0x25, 0x1E, 0x01, 0x76, 0x1B,
	0x08, 0x24, 0x27, 0x13, 0x54, 0x23, 0x2B, 0x28, 0x0C, 0x5C, 0x2E, 0x28,
	0x02, 0x28, 0x55, 0x22, 0x3C, 0x09, 0x2E, 0x22, 0x52, 0x08, 0x5B, 0x69,
	0x3A, 0x0B, 0x38, 0x2F, 0x73, 0x0F, 0x22, 0x57, 0x04, 0x15, 0x05, 0x59,
	0x24, 0x05, 0x13, 0x3F, 0x2C, 0x1F, 0x5B, 0x07, 0x25, 0x50, 0x09, 0x31,
	0x2F, 0x3D, 0x08, 0x28, 0x0D, 0x71, 0x0B, 0x11, 0x41, 0x00, 0x08, 0x3D,
	0x30, 0x19, 0x5B, 0x01, 0x1B, 0x29, 0x5F, 0x1D, 0x77, 0x28, 0x16, 0x5A,
	0x0D, 0x33, 0x0B, 0x2F, 0x09, 0x0E, 0x0E, 0x54, 0x24, 0x5E, 0x26, 0x08,
	0x36, 0x3B, 0x5D, 0x28, 0x3B, 0x5E, 0x59, 0x19, 0x3D, 0x30, 0x1D, 0x2D,
	0x39, 0x24, 0x2E, 0x1D, 0x23, 0x29, 0x05, 0x0A, 0x19, 0x2F, 0x08, 0x01,
	0x35, 0x1C, 0x2E, 0x18, 0x1B, 0x2F, 0x2A, 0x28, 0x0C, 0x26, 0x1A, 0x25,
	0x38, 0x3A, 0x1B, 0x76, 0x0F, 0x00, 0x0A, 0x3D, 0x21, 0x36, 0x35, 0x58,
	0x0F, 0x2A, 0x1C, 0x14, 0x58, 0x53, 0x05, 0x3C, 0x14, 0x39, 0x06, 0x08,
	0x5B, 0x2C, 0x0A, 0x23, 0x23, 0x09, 0x08, 0x04, 0x05, 0x3B, 0x04, 0x34,
	0x02, 0x24, 0x2F, 0x29, 0x39, 0x07, 0x26, 0x24, 0x2D, 0x14, 0x58, 0x0A,
	0x18, 0x1D, 0x38, 0x5A, 0x01, 0x11, 0x0A, 0x2D, 0x1F, 0x29, 0x15, 0x3A,
	0x54, 0x0F, 0x5D, 0x0A, 0x5F, 0x31, 0x1A, 0x2D, 0x23, 0x1D, 0x26, 0x28,
	0x25, 0x24, 0x3A, 0x27, 0x5C, 0x05, 0x09, 0x3F, 0x26, 0x1F, 0x5C, 0x2E,
	0x58, 0x07, 0x1E, 0x32, 0x14, 0x47, 0x17, 0x00, 0x22, 0x70, 0x03, 0x04,
	0x29, 0x1B, 0x3B, 0x27, 0x25, 0x3F, 0x06, 0x7B, 0x24, 0x13, 0x5E, 0x25,
	0x11, 0x1C, 0x33, 0x2A, 0x2C, 0x74, 0x58, 0x54, 0x38, 0x3B, 0x32, 0x26,
	0x30, 0x20, 0x28, 0x09, 0x5D, 0x34, 0x2F, 0x53, 0x0B, 0x43, 0x2C, 0x06,
	0x2F, 0x24, 0x0F, 0x57, 0x06, 0x3D, 0x76, 0x27, 0x25, 0x07, 0x38, 0x13,
	0x24, 0x08, 0x0D, 0x3B, 0x25, 0x29, 0x0B, 0x2D, 0x0C, 0x30, 0x5F, 0x11,
	0x0C, 0x3F, 0x71, 0x5F, 0x2F, 0x57, 0x1B, 0x31, 0x58, 0x20, 0x06, 0x1F,
	0x35, 0x47, 0x36, 0x38, 0x1D, 0x2D, 0x5F, 0x52, 0x1C, 0x05, 0x30, 0x03,
	0x07, 0x07, 0x02, 0x77, 0x2D, 0x39, 0x09, 0x12, 0x17, 0x59, 0x10, 0x37,
	0x2D, 0x23, 0x5F, 0x53, 0x19, 0x2E, 0x2B, 0x5B, 0x4E, 0x5B, 0x27, 0x75,
	0x22, 0x30, 0x26, 0x1D, 0x01, 0x0B, 0x57, 0x1D, 0x40, 0x0D, 0x1A, 0x17,
	0x00, 0x33, 0x2A, 0x16, 0x34, 0x05, 0x1E, 0x10, 0x1C, 0x04, 0x3D, 0x5A,
	0x38, 0x05, 0x02, 0x3B, 0x1D, 0x12, 0x00, 0x37, 0x41, 0x24, 0x0E, 0x2E,
	0x07, 0x17, 0x07, 0x09, 0x25, 0x13, 0x22, 0x0D, 0x21, 0x2E, 0x57, 0x1F,
	0x44, 0x25, 0x47, 0x28, 0x5D, 0x18, 0x38, 0x0A, 0x4E, 0x1A, 0x39, 0x3A,
	0x3D, 0x32, 0x29, 0x12, 0x38, 0x19, 0x07, 0x3D, 0x06, 0x23, 0x2F, 0x3B,
	0x14, 0x1C, 0x75, 0x06, 0x29, 0x23, 0x0F, 0x2D, 0x5D, 0x30, 0x03, 0x11,
	0x27, 0x19, 0x25, 0x21, 0x0D, 0x27, 0x3A, 0x56, 0x01, 0x39, 0x00, 0x0B,
	0x11, 0x29, 0x27, 0x23, 0x54, 0x0B, 0x01, 0x1B, 0x26, 0x43, 0x51, 0x3B,
	0x0D, 0x31, 0x02, 0x13, 0x28, 0x2C, 0x0D, 0x3C, 0x39, 0x5D, 0x59, 0x72,
	0x59, 0x33, 0x23, 0x3D, 0x0D, 0x2D, 0x02, 0x04, 0x0D, 0x31, 0x24, 0x18,
	0x0F, 0x3C, 0x72, 0x59, 0x0D, 0x45, 0x2A, 0x10, 0x3A, 0x12, 0x03, 0x12,
	0x71, 0x5A, 0x0C, 0x5E, 0x3B, 0x75, 0x1C, 0x2E, 0x45, 0x5E, 0x04, 0x59,
	0x22, 0x57, 0x5C, 0x01, 0x28, 0x54, 0x1E, 0x18, 0x74, 0x01, 0x35, 0x21,
	0x5E, 0x76, 0x2F, 0x26, 0x28, 0x3B, 0x35, 0x19, 0x18, 0x02, 0x52, 0x28,
	0x55, 0x11, 0x1A, 0x27, 0x06, 0x05, 0x57, 0x09, 0x25, 0x26, 0x14, 0x24,
	0x23, 0x0D, 0x24, 0x1D, 0x28, 0x3C, 0x44, 0x1B, 0x19, 0x29, 0x27, 0x2D,
	0x33, 0x0A, 0x08, 0x5F, 0x58, 0x10, 0x24, 0x10, 0x2B, 0x5B, 0x01, 0x07,
	0x54, 0x06, 0x33, 0x00, 0x43, 0x2A, 0x5D, 0x27, 0x31, 0x5A, 0x08, 0x05,
	0x23, 0x7A, 0x00, 0x12, 0x1F, 0x40, 0x2A, 0x1D, 0x18, 0x0F, 0x27, 0x30,
	0x5D, 0x12, 0x59, 0x53, 0x03, 0x3B, 0x35, 0x3D, 0x44, 0x01, 0x5B, 0x08,
	0x45, 0x1F, 0x00, 0x34, 0x0A, 0x20, 0x26, 0x20, 0x0D, 0x4A, 0x0F, 0x03,
	0x2C, 0x38, 0x11, 0x57, 0x2A, 0x15, 0x5C, 0x26, 0x24, 0x1B, 0x0A, 0x06,
	0x10, 0x3D, 0x1B, 0x2D, 0x1C, 0x24, 0x56, 0x5F, 0x72, 0x1C, 0x34, 0x0C,
	0x0F, 0x0D, 0x2A, 0x33, 0x1C, 0x1D, 0x0D, 0x1B, 0x2A, 0x2A, 0x1E, 0x16,
	0x1A, 0x51, 0x45, 0x40, 0x01, 0x20, 0x0B, 0x1E, 0x01, 0x3A, 0x1F, 0x52,
	0x1D, 0x23, 0x7A, 0x03, 0x4A, 0x2C, 0x44, 0x3A, 0x35, 0x3B, 0x09, 0x2A,
	0x05, 0x54, 0x2D, 0x27, 0x5C, 0x32, 0x16, 0x36, 0x22, 0x5A, 0x77, 0x43,
	0x28, 0x41, 0x1F, 0x28, 0x47, 0x12, 0x39, 0x09, 0x10, 0x08, 0x30, 0x34,
	0x5A, 0x0D, 0x54, 0x31, 0x22, 0x40, 0x0C, 0x26, 0x58, 0x25, 0x3B, 0x17,
	0x1C, 0x53, 0x58, 0x5C, 0x70, 0x1A, 0x20, 0x3A, 0x28, 0x28, 0x1E, 0x0B,
	0x1F, 0x23, 0x2E, 0x5A, 0x15, 0x06, 0x44, 0x32, 0x5C, 0x36, 0x1A, 0x2F,
	0x1B, 0x3C, 0x14, 0x56, 0x25, 0x03, 0x16, 0x29, 0x3F, 0x29, 0x38, 0x2F,
	0x2C, 0x3B, 0x07, 0x15, 0x14, 0x33, 0x23, 0x2F, 0x17, 0x16, 0x03, 0x1E,
	0x24, 0x0A, 0x0D, 0x50, 0x3C, 0x3D, 0x70, 0x14, 0x34, 0x3D, 0x1C, 0x77,
	0x08, 0x07, 0x59, 0x5C, 0x1A, 0x39, 0x24, 0x06, 0x04, 0x72, 0x3C, 0x25,
	0x2D, 0x1A, 0x3A, 0x25, 0x52, 0x21, 0x02, 0x34, 0x28, 0x0E, 0x57, 0x0E,
	0x29, 0x03, 0x59, 0x1F, 0x1A, 0x18, 0x09, 0x58, 0x07, 0x0D, 0x04, 0x01,
	0x51, 0x2C, 0x44, 0x33, 0x5D, 0x2C, 0x3E, 0x5A, 0x3B, 0x2F, 0x54, 0x18,
	0x29, 0x11, 0x28, 0x28, 0x00, 0x18, 0x27, 0x35, 0x28, 0x5D, 0x23, 0x27,
	0x3B, 0x4A, 0x04, 0x5D, 0x71, 0x3A, 0x15, 0x27, 0x24, 0x76, 0x06, 0x3B,
	0x27, 0x08, 0x2F, 0x0E, 0x51, 0x16, 0x40, 0x05, 0x06, 0x04, 0x34, 0x2C,
	0x10, 0x01, 0x20, 0x24, 0x00, 0x29, 0x29, 0x11, 0x1D, 0x02, 0x37, 0x54,
	0x37, 0x5C, 0x01, 0x08, 0x23, 0x1B, 0x07, 0x3F, 0x1B, 0x15, 0x4A, 0x3C,
	0x19, 0x0E, 0x16, 0x50, 0x22, 0x3F, 0x73, 0x55, 0x3B, 0x56, 0x31, 0x2F,
	0x3B, 0x37, 0x20, 0x53, 0x07, 0x5D, 0x06, 0x21, 0x1C, 0x7B, 0x43, 0x22,
	0x3F, 0x12, 0x6D, 0x55, 0x25, 0x5A, 0x2A, 0x27, 0x5C, 0x50, 0x17, 0x1E,
	0x07, 0x5C, 0x4E, 0x3B, 0x02, 0x29, 0x25, 0x09, 0x21, 0x0C, 0x31, 0x0F,
	0x26, 0x2F, 0x20, 0x00, 0x09, 0x2A, 0x3B, 0x3F, 0x71, 0x2F, 0x20, 0x08,
	0x24, 0x04, 0x09, 0x2D, 0x5D, 0x1D, 0x29, 0x00, 0x50, 0x2C, 0x0E, 0x25,
	0x3C, 0x26, 0x58, 0x04, 0x13, 0x3E, 0x2E, 0x04, 0x5E, 0x12, 0x58, 0x15,
	0x05, 0x26, 0x08, 0x38, 0x08, 0x5B, 0x33, 0x1B, 0x35, 0x15, 0x29, 0x33,
	0x0C, 0x07, 0x15, 0x02, 0x26, 0x26, 0x59, 0x1B, 0x1E, 0x19, 0x74, 0x26,
	0x2B, 0x05, 0x02, 0x0E, 0x59, 0x25, 0x36, 0x3A, 0x69, 0x36, 0x11, 0x3C,
	0x58, 0x33, 0x38, 0x36, 0x59, 0x2D, 0x33, 0x5D, 0x05, 0x3C, 0x3E, 0x0B,
	0x39, 0x1B, 0x03, 0x1D, 0x75, 0x07, 0x52, 0x3B, 0x24, 0x12, 0x0E, 0x08,
	0x24, 0x18, 0x06, 0x2D, 0x02, 0x45, 0x09, 0x16, 0x0E, 0x59, 0x26, 0x11,
	0x20, 0x3D, 0x2B, 0x21, 0x08, 0x11, 0x47, 0x2C, 0x3B, 0x18, 0x29, 0x0E,
	0x0D, 0x37, 0x53, 0x0A, 0x02, 0x0D, 0x0A, 0x5C, 0x13, 0x07, 0x54, 0x0D,
	0x2F, 0x31, 0x08, 0x19, 0x39, 0x22, 0x76, 0x06, 0x03, 0x45, 0x26, 0x29,
	0x21, 0x0D, 0x57, 0x28, 0x09, 0x1F, 0x0F, 0x3C, 0x22, 0x3A, 0x1C, 0x56,
	0x56, 0x5C, 0x20, 0x3C, 0x33, 0x37, 0x1D, 0x76, 0x1D, 0x2E, 0x3A, 0x52,
	0x01, 0x1F, 0x0A, 0x03, 0x31, 0x0E, 0x1E, 0x0E, 0x24, 0x0D, 0x1B, 0x55,
	0x2F, 0x1B, 0x3D, 0x7A, 0x14, 0x2E, 0x00, 0x00, 0x76, 0x2E, 0x37, 0x06,
	0x3B, 0x29, 0x43, 0x51, 0x2F, 0x1E, 0x30, 0x07, 0x12, 0x17, 0x06, 0x21,
	0x58, 0x18, 0x09, 0x53, 0x72, 0x06, 0x0F, 0x00, 0x0C, 0x1B, 0x26, 0x09,
	0x57, 0x12, 0x21, 0x5A, 0x58, 0x07, 0x21, 0x15, 0x20, 0x24, 0x28, 0x27,
	0x25, 0x22, 0x29, 0x2C, 0x2F, 0x2C, 0x35, 0x4A, 0x01, 0x01, 0x0E, 0x3E,
	0x3B, 0x04, 0x05, 0x28, 0x34, 0x22, 0x0C, 0x03, 0x31, 0x0D, 0x0F, 0x1B,
	0x0C, 0x03, 0x2A, 0x2A, 0x58, 0x00, 0x21, 0x20, 0x0C, 0x27, 0x08, 0x3A,
	0x5E, 0x20, 0x3B, 0x1C, 0x27, 0x09, 0x32, 0x57, 0x0A, 0x12, 0x1D, 0x0D,
	0x21, 0x00, 0x03, 0x02, 0x34, 0x3E, 0x20, 0x27, 0x0A, 0x51, 0x3E, 0x09,
	0x3B, 0x54, 0x0D, 0x2B, 0x52, 0x71, 0x2D, 0x0D, 0x36, 0x44, 0x1B, 0x0F,
	0x02, 0x14, 0x11, 0x25, 0x00, 0x0C, 0x3B, 0x19, 0x37, 0x3F, 0x2D, 0x29,
	0x1D, 0x74, 0x29, 0x27, 0x3E, 0x3D, 0x20, 0x15, 0x09, 0x39, 0x53, 0x35,
	0x1F, 0x18, 0x34, 0x5C, 0x27, 0x14, 0x25, 0x3B, 0x07, 0x21, 0x0F, 0x23,
	0x41, 0x40, 0x70, 0x00, 0x57, 0x09, 0x25, 0x20, 0x5E, 0x2A, 0x37, 0x1B,
	0x01, 0x04, 0x33, 0x36, 0x1E, 0x13, 0x5A, 0x0D, 0x06, 0x06, 0x0D, 0x5F,
	0x16, 0x03, 0x08, 0x34, 0x35, 0x2D, 0x14, 0x5F, 0x06, 0x09, 0x09, 0x3D,
	0x3F, 0x2C, 0x5C, 0x2E, 0x03, 0x07, 0x14, 0x34, 0x0F, 0x1F, 0x21, 0x13,
	0x07, 0x2B, 0x22, 0x3D, 0x11, 0x2A, 0x0B, 0x16, 0x44, 0x25, 0x1A, 0x20,
	0x1E, 0x0C, 0x0B, 0x00, 0x59, 0x56, 0x11, 0x30, 0x5E, 0x0E, 0x34, 0x5B,
	0x2C, 0x15, 0x56, 0x01, 0x5B, 0x0E, 0x16, 0x26, 0x24, 0x07, 0x69, 0x0A,
	0x2A, 0x23, 0x00, 0x77, 0x0E, 0x18, 0x1E, 0x5D, 0x30, 0x1C, 0x28, 0x3F,
	0x03, 0x70, 0x15, 0x10, 0x38, 0x3C, 0x26, 0x35, 0x31, 0x24, 0x3F, 0x01,
	0x3B, 0x58, 0x56, 0x22, 0x0D, 0x1B, 0x15, 0x19, 0x26, 0x1A, 0x29, 0x37,
	0x56, 0x31, 0x77, 0x5F, 0x32, 0x2F, 0x11, 0x17, 0x1F, 0x19, 0x5C, 0x13,
	0x2A, 0x0D, 0x4E, 0x01, 0x53, 0x20, 0x5A, 0x37, 0x5F, 0x5A, 0x05, 0x14,
	0x11, 0x21, 0x53, 0x16, 0x1A, 0x31, 0x09, 0x20, 0x7A, 0x5A, 0x28, 0x23,
	0x0C, 0x76, 0x01, 0x0E, 0x28, 0x5C, 0x0C, 0x25, 0x10, 0x0A, 0x06, 0x34,
	0x21, 0x19, 0x0B, 0x24, 0x18, 0x58, 0x38, 0x1B, 0x23, 0x06, 0x3E, 0x54,
	0x29, 0x13, 0x77, 0x21, 0x22, 0x41, 0x2C, 0x01, 0x19, 0x18, 0x1B, 0x27,
	0x2C, 0x05, 0x16, 0x59, 0x29, 0x2F, 0x18, 0x55, 0x17, 0x3D, 0x37, 0x58,
	0x09, 0x09, 0x40, 0x6D, 0x2F, 0x26, 0x25, 0x19, 0x2B, 0x09, 0x2A, 0x2A,
	0x3F, 0x1A, 0x5D, 0x07, 0x5E, 0x09, 0x23, 0x2D, 0x35, 0x1A, 0x28, 0x2A,
	0x3B, 0x0D, 0x3E, 0x59, 0x74, 0x5E, 0x19, 0x3A, 0x11, 0x71, 0x5C, 0x04,
	0x20, 0x22, 0x6D, 0x5D, 0x31, 0x38, 0x44, 0x3B, 0x14, 0x28, 0x2D, 0x1E,
	0x1A, 0x29, 0x20, 0x36, 0x33, 0x25, 0x08, 0x28, 0x16, 0x01, 0x37, 0x38,
	0x57, 0x0F, 0x27, 0x74, 0x2F, 0x00, 0x39, 0x38, 0x7B, 0x43, 0x26, 0x5B,
	0x04, 0x28, 0x0A, 0x50, 0x56, 0x1F, 0x24, 0x28, 0x0C, 0x45, 0x08, 0x00,
	0x04, 0x38, 0x18, 0x12, 0x16, 0x5C, 0x0F, 0x16, 0x2E, 0x33, 0x29, 0x0D,
	0x5B, 0x2C, 0x3A, 0x1E, 0x35, 0x37, 0x28, 0x71, 0x20, 0x13, 0x04, 0x3D,
	0x2B, 0x1C, 0x04, 0x5D, 0x02, 0x7B, 0x25, 0x16, 0x3E, 0x1B, 0x16, 0x24,
	0x02, 0x5A, 0x5C, 0x2A, 0x2F, 0x0F, 0x56, 0x53, 0x16, 0x5B, 0x14, 0x17,
	0x5E, 0x17, 0x2D, 0x04, 0x08, 0x31, 0x06, 0x02, 0x14, 0x3B, 0x18, 0x29,
	0x19, 0x0F, 0x0C, 0x07, 0x33, 0x5A, 0x2E, 0x27, 0x1A, 0x2C, 0x14, 0x58,
	0x26, 0x03, 0x75, 0x1A, 0x59, 0x5E, 0x12, 0x04, 0x08, 0x15, 0x3D, 0x58,
	0x04, 0x5E, 0x2F, 0x56, 0x2F, 0x75, 0x39, 0x11, 0x25, 0x31, 0x10, 0x29,
	0x28, 0x17, 0x11, 0x07, 0x2B, 0x29, 0x5C, 0x33, 0x1A, 0x15, 0x02, 0x20,
	0x26, 0x75, 0x58, 0x2C, 0x2F, 0x13, 0x0A, 0x0F, 0x12, 0x17, 0x05, 0x11,
	0x15, 0x35, 0x3A, 0x03, 0x0C, 0x0F, 0x33, 0x21, 0x3D, 0x2A, 0x15, 0x34,
	0x3A, 0x3B, 0x7B, 0x47, 0x30, 0x5A, 0x39, 0x6D, 0x54, 0x1B, 0x37, 0x32,
	0x29, 0x2A, 0x09, 0x34, 0x3C, 0x0B, 0x1C, 0x55, 0x1B, 0x5F, 0x09, 0x26,
	0x28, 0x25, 0x26, 0x1A, 0x19, 0x09, 0x24, 0x5A, 0x16, 0x3E, 0x2A, 0x17,
	0x2A, 0x35, 0x39, 0x34, 0x04, 0x18, 0x24, 0x1B, 0x39, 0x23, 0x3A, 0x06,
	0x0D, 0x36, 0x34, 0x19, 0x33, 0x2E, 0x03, 0x3C, 0x32, 0x03, 0x05, 0x33,
	0x08, 0x3C, 0x07, 0x1C, 0x58, 0x36, 0x00, 0x77, 0x1F, 0x0B, 0x59, 0x5D,
	0x70, 0x1C, 0x2D, 0x09, 0x40, 0x1B, 0x3E, 0x50, 0x5F, 0x1C, 0x3B, 0x29,
	0x27, 0x3E, 0x1C, 0x2D, 0x36, 0x2D, 0x01, 0x26, 0x35, 0x27, 0x17, 0x23,
	0x1B, 0x7A, 0x55, 0x20, 0x29, 0x1A, 0x69, 0x08, 0x1B, 0x00, 0x26, 0x18,
	0x5D, 0x38, 0x1C, 0x1B, 0x33, 0x19, 0x0D, 0x27, 0x3F, 0x70, 0x3B, 0x16,
	0x3C, 0x23, 0x0F, 0x54, 0x04, 0x2C, 0x5A, 0x14, 0x5A, 0x4A, 0x56, 0x21,
	0x05, 0x25, 0x1B, 0x5D, 0x0F, 0x03, 0x20, 0x56, 0x5C, 0x26, 0x3A, 0x16,
	0x37, 0x05, 0x1E, 0x18, 0x3A, 0x03, 0x07, 0x59, 0x06, 0x24, 0x08, 0x59,
	0x19, 0x31, 0x03, 0x56, 0x3D, 0x1B, 0x26, 0x08, 0x2A, 0x41, 0x26, 0x7B,
	0x03, 0x2C, 0x1F, 0x21, 0x2D, 0x5B, 0x28, 0x16, 0x25, 0x0B, 0x5F, 0x0F,
	0x2D, 0x1E, 0x10, 0x0D, 0x54, 0x27, 0x04, 0x03, 0x29, 0x00, 0x18, 0x18,
	0x14, 0x16, 0x4E, 0x45, 0x22, 0x2A, 0x3E, 0x08, 0x07, 0x5A, 0x38, 0x21,
	0x05, 0x06, 0x1B, 0x12, 0x1A, 0x57, 0x34, 0x5E, 0x2A, 0x01, 0x20, 0x1E,
	0x2D, 0x31, 0x5F, 0x4E, 0x39, 0x53, 0x69, 0x3D, 0x53, 0x25, 0x5A, 0x12,
	0x09, 0x38, 0x2C, 0x1E, 0x0C, 0x2A, 0x39, 0x5A, 0x5C, 0x69, 0x0D, 0x35,
	0x1D, 0x58, 0x0A, 0x15, 0x07, 0x2A, 0x19, 0x05, 0x0F, 0x16, 0x5A, 0x04,
	0x09, 0x15, 0x2D, 0x3E, 0x33, 0x0B, 0x58, 0x18, 0x36, 0x38, 0x3A, 0x2E,
	0x26, 0x19, 0x11, 0x26, 0x03, 0x04, 0x23, 0x25, 0x16, 0x38, 0x0E, 0x58,
	0x5B, 0x0B, 0x2A, 0x52, 0x26, 0x1A, 0x2D, 0x34, 0x30, 0x0B, 0x53, 0x00,
	0x5D, 0x19, 0x05, 0x25, 0x7B, 0x02, 0x38, 0x2A, 0x2D, 0x6D, 0x5F, 0x02,
	0x04, 0x52, 0x26, 0x58, 0x03, 0x29, 0x04, 0x01, 0x1C, 0x59, 0x58, 0x23,
	0x31, 0x09, 0x23, 0x39, 0x04, 0x15, 0x26, 0x2A, 0x09, 0x22, 0x05, 0x26,
	0x2B, 0x36, 0x05, 0x21, 0x5D, 0x35, 0x16, 0x0F, 0x75, 0x01, 0x2C, 0x38,
	0x5E, 0x33, 0x54, 0x14, 0x5F, 0x24, 0x71, 0x2A, 0x14, 0x58, 0x3B, 0x21,
	0x22, 0x59, 0x23, 0x32, 0x31, 0x1A, 0x27, 0x19, 0x06, 0x10, 0x34, 0x51,
	0x5D, 0x12, 0x30, 0x39, 0x07, 0x59, 0x58, 0x05, 0x1A, 0x02, 0x21, 0x3A,
	0x73, 0x5E, 0x4A, 0x3A, 0x5E, 0x03, 0x2E, 0x4A, 0x17, 0x59, 0x0B, 0x5F,
	0x2A, 0x22, 0x44, 0x2F, 0x07, 0x26, 0x00, 0x52, 0x12, 0x26, 0x54, 0x1B,
	0x3C, 0x30, 0x01, 0x38, 0x0C, 0x3A, 0x73, 0x55, 0x25, 0x0F, 0x3B, 0x73,
	0x34, 0x10, 0x08, 0x2F, 0x71, 0x34, 0x52, 0x3F, 0x1E, 0x73, 0x5C, 0x2D,
	0x23, 0x31, 0x15, 0x08, 0x32, 0x24, 0x5C, 0x21, 0x0B, 0x0B, 0x07, 0x3C,
	0x06, 0x0B, 0x38, 0x0C, 0x29, 0x28, 0x25, 0x55, 0x28, 0x5B, 0x2F, 0x5A,
	0x0E, 0x23, 0x58, 0x3B, 0x0D, 0x52, 0x2B, 0x1F, 0x0C, 0x2D, 0x02, 0x0D,
	0x1A, 0x6D, 0x3E, 0x37, 0x5D, 0x25, 0x04, 0x3D, 0x0C, 0x37, 0x3B, 0x26,
	0x2A, 0x16, 0x5A, 0x0A, 0x33, 0x01, 0x25, 0x45, 0x52, 0x18, 0x00, 0x12,
	0x3E, 0x5D, 0x03, 0x43, 0x2E, 0x57, 0x0E, 0x17, 0x05, 0x06, 0x18, 0x31,
	0x08, 0x5B, 0x2D, 0x41, 0x1A, 0x70, 0x3B, 0x26, 0x57, 0x21, 0x0A, 0x22,
	0x2B, 0x14, 0x3D, 0x37, 0x59, 0x18, 0x02, 0x18, 0x77, 0x2F, 0x02, 0x3D,
	0x2C, 0x29, 0x1B, 0x50, 0x1D, 0x5D, 0x34, 0x1C, 0x59, 0x2A, 0x5F, 0x28,
	0x01, 0x4E, 0x57, 0x22, 0x29, 0x0B, 0x30, 0x5C, 0x59, 0x01, 0x3B, 0x14,
	0x18, 0x28, 0x15, 0x3A, 0x11, 0x21, 0x22, 0x24, 0x0B, 0x27, 0x03, 0x59,
	0x1A, 0x0F, 0x37, 0x14, 0x0D, 0x1A, 0x5D, 0x08, 0x16, 0x19, 0x30, 0x25,
	0x27, 0x28, 0x3E, 0x34, 0x01, 0x4A, 0x27, 0x1D, 0x14, 0x23, 0x07, 0x5D,
	0x21, 0x0E, 0x1A, 0x14, 0x2A, 0x2A, 0x35, 0x0D, 0x23, 0x07, 0x44, 0x0F,
	0x1B, 0x14, 0x56, 0x23, 0x13, 0x3E, 0x2E, 0x2D, 0x38, 0x72, 0x0F, 0x29,
	0x3A, 0x39, 0x69, 0x3C, 0x2F, 0x1C, 0x24, 0x31, 0x3D, 0x1B, 0x3E, 0x1D,
	0x31, 0x5E, 0x38, 0x56, 0x3C, 0x69, 0x0B, 0x20, 0x58, 0x21, 0x73, 0x16,
	0x0C, 0x0C, 0x44, 0x34, 0x21, 0x2A, 0x00, 0x59, 0x16, 0x5F, 0x50, 0x29,
	0x33, 0x01, 0x2D, 0x07, 0x5D, 0x1F, 0x11, 0x2E, 0x13, 0x5C, 0x3B, 0x69,
	0x43, 0x30, 0x1E, 0x1C, 0x25, 0x0F, 0x4E, 0x0C, 0x5F, 0x31, 0x54, 0x13,
	0x26, 0x00, 0x76, 0x3F, 0x52, 0x20, 0x44, 0x25, 0x15, 0x15, 0x3C, 0x06,
	0x69, 0x54, 0x25, 0x0B, 0x52, 0x28, 0x0F, 0x0C, 0x5C, 0x0E, 0x1A, 0x06,
	0x2F, 0x03, 0x52, 0x11, 0x09, 0x19, 0x56, 0x3B, 0x0A, 0x39, 0x10, 0x38,
	0x1E, 0x30, 0x5D, 0x05, 0x04, 0x01, 0x05, 0x09, 0x52, 0x06, 0x2E, 0x74,
	0x07, 0x37, 0x5E, 0x1C, 0x37, 0x07, 0x0A, 0x04, 0x1C, 0x3A, 0x5A, 0x17,
	0x37, 0x1E, 0x38, 0x0B, 0x51, 0x58, 0x0E, 0x18, 0x07, 0x27, 0x36, 0x12,
	0x7B, 0x1E, 0x16, 0x3D, 0x2F, 0x32, 0x16, 0x1B, 0x29, 0x02, 0x69, 0x5A,
	0x22, 0x1D, 0x0D, 0x14, 0x14, 0x18, 0x57, 0x0A, 0x73, 0x0B, 0x0F, 0x1B,
	0x2D, 0x23, 0x09, 0x33, 0x2D, 0x52, 0x2C, 0x02, 0x53, 0x18, 0x2F, 0x0B,
	0x5A, 0x39, 0x29, 0x5C, 0x2D, 0x1E, 0x04, 0x5B, 0x12, 0x2D, 0x2E, 0x07,
	0x14, 0x00, 0x24, 0x0D, 0x29, 0x1B, 0x5B, 0x26, 0x01, 0x10, 0x04, 0x0F,
	0x03, 0x58, 0x07, 0x36, 0x53, 0x6D, 0x02, 0x15, 0x56, 0x0C, 0x29, 0x18,
	0x36, 0x20, 0x0D, 0x2F, 0x3C, 0x58, 0x2C, 0x09, 0x32, 0x2F, 0x53, 0x0C,
	0x58, 0x10, 0x3F, 0x0E, 0x39, 0x44, 0x24, 0x5B, 0x58, 0x0A, 0x5A, 0x69,
	0x1D, 0x2C, 0x21, 0x03, 0x70, 0x2B, 0x20, 0x3F, 0x25, 0x18, 0x26, 0x22,
	0x57, 0x33, 0x07, 0x5F, 0x3B, 0x2A, 0x23, 0x27, 0x09, 0x2C, 0x1C, 0x22,
	0x73, 0x24, 0x52, 0x59, 0x5D, 0x13, 0x06, 0x52, 0x2D, 0x2C, 0x35, 0x29,
	0x17, 0x02, 0x00, 0x16, 0x1D, 0x25, 0x05, 0x3A, 0x2F, 0x24, 0x26, 0x0F,
	0x2E, 0x0C, 0x01, 0x3B, 0x28, 0x04, 0x12, 0x29, 0x0C, 0x34, 0x26, 0x00,
	0x05, 0x00, 0x1B, 0x33, 0x74, 0x3A, 0x23, 0x0B, 0x24, 0x08, 0x55, 0x0C,
	0x19, 0x02, 0x16, 0x0B, 0x30, 0x16, 0x05, 0x2E, 0x38, 0x04, 0x5E, 0x5A,
	0x0D, 0x39, 0x29, 0x2A, 0x0F, 0x7B, 0x1E, 0x50, 0x38, 0x5C, 0x2B, 0x36,
	0x18, 0x24, 0x0E, 0x25, 0x0E, 0x2C, 0x19, 0x58, 0x30, 0x55, 0x33, 0x36,
	0x3C, 0x14, 0x5F, 0x2D, 0x5E, 0x13, 0x04, 0x2E, 0x54, 0x24, 0x5D, 0x01,
	0x0F, 0x3B, 0x3C, 0x24, 0x0D, 0x1F, 0x10, 0x2D, 0x03, 0x74, 0x0A, 0x2D,
	0x09, 0x19, 0x03, 0x23, 0x17, 0x17, 0x5F, 0x2B, 0x21, 0x11, 0x14, 0x03,
	0x13, 0x0F, 0x18, 0x56, 0x29, 0x33, 0x3F, 0x24, 0x2F, 0x58, 0x76, 0x1C,
	0x10, 0x3D, 0x1F, 0x24, 0x3D, 0x17, 0x41, 0x27, 0x36, 0x35, 0x0A, 0x2C,
	0x52, 0x35, 0x01, 0x59, 0x0C, 0x3B, 0x72, 0x55, 0x2D, 0x5B, 0x2D, 0x2C,
	0x54, 0x12, 0x18, 0x00, 0x15, 0x19, 0x09, 0x59, 0x3E, 0x0B, 0x0A, 0x02,
	0x3B, 0x05, 0x72, 0x0A, 0x57, 0x09, 0x09, 0x69, 0x0D, 0x20, 0x03, 0x2D,
	0x09, 0x3C, 0x03, 0x09, 0x2D, 0x09, 0x3F, 0x10, 0x56, 0x11, 0x03, 0x26,
	0x25, 0x14, 0x3F, 0x25, 0x1B, 0x36, 0x27, 0x0A, 0x2D, 0x08, 0x07, 0x5A,
	0x05, 0x38, 0x47, 0x33, 0x2C, 0x39, 0x0B, 0x58, 0x50, 0x2A, 0x09, 0x7A,
	0x5A, 0x28, 0x09, 0x19, 0x75, 0x58, 0x0C, 0x36, 0x5D, 0x26, 0x2D, 0x09,
	0x1E, 0x3A, 0x2F, 0x09, 0x13, 0x28, 0x32, 0x0F, 0x0D, 0x4E, 0x2B, 0x29,
	0x2D, 0x5F, 0x50, 0x16, 0x20, 0x29, 0x54, 0x0B, 0x5D, 0x3A, 0x2B, 0x22,
	0x23, 0x1A, 0x0A, 0x24, 0x1C, 0x31, 0x20, 0x3F, 0x0F, 0x3C, 0x4A, 0x1E,
	0x5F, 0x24, 0x01, 0x52, 0x1D, 0x2D, 0x71, 0x28, 0x15, 0x1A, 0x26, 0x1B,
	0x25, 0x27, 0x5F, 0x21, 0x21, 0x2D, 0x07, 0x5E, 0x2D, 0x2E, 0x5D, 0x35,
	0x5E, 0x1C, 0x05, 0x5E, 0x3B, 0x45, 0x25, 0x0C, 0x09, 0x30, 0x16, 0x11,
	0x03, 0x1B, 0x39, 0x5A, 0x1E, 0x70, 0x3D, 0x2F, 0x07, 0x5D, 0x2D, 0x23,
	0x23, 0x26, 0x27, 0x0D, 0x25, 0x2D, 0x34, 0x1F, 0x2E, 0x2D, 0x0A, 0x0C,
	0x58, 0x35, 0x1B, 0x32, 0x20, 0x1E, 0x75, 0x59, 0x09, 0x28, 0x2F, 0x2A,
	0x0A, 0x16, 0x07, 0x2D, 0x73, 0x5D, 0x4E, 0x28, 0x44, 0x04, 0x43, 0x0C,
	0x2F, 0x2F, 0x18, 0x15, 0x3B, 0x19, 0x01, 0x05, 0x05, 0x19, 0x5C, 0x0F,
	0x35, 0x28, 0x09, 0x5D, 0x0A, 0x16, 0x15, 0x2C, 0x1D, 0x40, 0x03, 0x55,
	0x59, 0x2C, 0x1A, 0x26, 0x22, 0x1B, 0x03, 0x20, 0x11, 0x27, 0x03, 0x45,
	0x52, 0x00, 0x5D, 0x4A, 0x20, 0x23, 0x07, 0x5A, 0x57, 0x3E, 0x38, 0x00,
	0x5C, 0x02, 0x5E, 0x18, 0x1A, 0x1C, 0x37, 0x1E, 0x40, 0x29, 0x1D, 0x10,
	0x21, 0x21, 0x24, 0x1C, 0x25, 0x06, 0x02, 0x2C, 0x2E, 0x0C, 0x1E, 0x2F,
	0x71, 0x00, 0x18, 0x03, 0x26, 0x0E, 0x04, 0x07, 0x1E, 0x33, 0x26, 0x38,
	0x55, 0x3B, 0x1F, 0x0F, 0x2E, 0x15, 0x27, 0x52, 0x37, 0x22, 0x57, 0x06,
	0x18, 0x32, 0x20, 0x57, 0x17, 0x03, 0x11, 0x09, 0x51, 0x14, 0x3D, 0x20,
	0x08, 0x0B, 0x59, 0x33, 0x08, 0x5F, 0x22, 0x00, 0x3B, 0x2B, 0x1E, 0x31,
	0x3F, 0x2F, 0x27, 0x1B, 0x56, 0x26, 0x39, 0x21, 0x02, 0x03, 0x5F, 0x3C,
	0x34, 0x3B, 0x16, 0x3A, 0x03, 0x14, 0x21, 0x02, 0x1A, 0x03, 0x3B, 0x0A,
	0x0F, 0x09, 0x05, 0x3B, 0x55, 0x4E, 0x23, 0x1B, 0x37, 0x20, 0x14, 0x5B,
	0x52, 0x30, 0x02, 0x0A, 0x05, 0x19, 0x38, 0x3A, 0x54, 0x3A, 0x04, 0x0D,
	0x1E, 0x34, 0x36, 0x29, 0x31, 0x58, 0x0C, 0x0A, 0x5D, 0x2C, 0x04, 0x30,
	0x06, 0x1F, 0x0A, 0x43, 0x54, 0x19, 0x44, 0x76, 0x0F, 0x4A, 0x09, 0x33,
	0x7B, 0x22, 0x2B, 0x0B, 0x28, 0x15, 0x39, 0x58, 0x5C, 0x59, 0x24, 0x5C,
	0x1B, 0x2A, 0x0C, 0x37, 0x16, 0x22, 0x00, 0x3C, 0x2D, 0x3B, 0x38, 0x16,
	0x08, 0x03, 0x1E, 0x31, 0x16, 0x33, 0x73, 0x0A, 0x32, 0x2D, 0x5A, 0x69,
	0x01, 0x54, 0x01, 0x44, 0x03, 0x23, 0x15, 0x0B, 0x1A, 0x2F, 0x0B, 0x2E,
	0x57, 0x2D, 0x34, 0x03, 0x4A, 0x20, 0x3C, 0x18, 0x15, 0x39, 0x3A, 0x13,
	0x15, 0x01, 0x4A, 0x28, 0x3B, 0x38, 0x29, 0x3B, 0x22, 0x11, 0x05, 0x16,
	0x30, 0x00, 0x0D, 0x01, 0x5F, 0x29, 0x26, 0x00, 0x14, 0x3F, 0x19, 0x5B,
	0x00, 0x27, 0x5D, 0x06, 0x14, 0x5F, 0x1B, 0x5F, 0x2F, 0x0B, 0x18, 0x16,
	0x5B, 0x30, 0x37, 0x2E, 0x05, 0x23, 0x51, 0x08, 0x12, 0x3B, 0x04, 0x24,
	0x57, 0x08, 0x7A, 0x34, 0x58, 0x36, 0x39, 0x38, 0x16, 0x57, 0x23, 0x39,
	0x27, 0x58, 0x09, 0x1A, 0x09, 0x2F, 0x34, 0x27, 0x00, 0x3A, 0x6D, 0x19,
	0x2A, 0x17, 0x1B, 0x09, 0x08, 0x2B, 0x20, 0x27, 0x72, 0x06, 0x00, 0x5B,
	0x18, 0x2E, 0x43, 0x24, 0x36, 0x08, 0x09, 0x0B, 0x1B, 0x01, 0x5D, 0x20,
	0x34, 0x2A, 0x23, 0x3E, 0x35, 0x43, 0x03, 0x19, 0x21, 0x32, 0x0A, 0x2F,
	0x0B, 0x58, 0x12, 0x25, 0x33, 0x1E, 0x1F, 0x21, 0x07, 0x0D, 0x2D, 0x1C,
	0x38, 0x0F, 0x55, 0x5C, 0x1E, 0x26, 0x59, 0x08, 0x03, 0x5A, 0x38, 0x0E,
	0x0F, 0x0B, 0x52, 0x17, 0x54, 0x12, 0x2B, 0x33, 0x2F, 0x0F, 0x3B, 0x38,
	0x12, 0x16, 0x0A, 0x20, 0x22, 0x5E, 0x74, 0x1C, 0x38, 0x0F, 0x18, 0x2B,
	0x05, 0x38, 0x23, 0x05, 0x2A, 0x16, 0x04, 0x23, 0x29, 0x29, 0x5D, 0x0C,
	0x00, 0x5A, 0x29, 0x1E, 0x18, 0x34, 0x1F, 0x18, 0x14, 0x0C, 0x2A, 0x04,
	0x34, 0x2E, 0x0B, 0x5B, 0x13, 0x10, 0x1B, 0x20, 0x5D, 0x3A, 0x17, 0x39,
	0x19, 0x45, 0x32, 0x21, 0x1C, 0x17, 0x2D, 0x2C, 0x3B, 0x35, 0x1B, 0x24,
	0x19, 0x21, 0x0A, 0x15, 0x3D, 0x3F, 0x76, 0x0E, 0x57, 0x57, 0x2F, 0x26,
	0x1B, 0x36, 0x2C, 0x58, 0x38, 0x1B, 0x3B, 0x22, 0x3B, 0x23, 0x55, 0x20,
	0x1F, 0x12, 0x34, 0x16, 0x4E, 0x3D, 0x2F, 0x12, 0x1F, 0x30, 0x1E, 0x0A,
	0x69, 0x23, 0x34, 0x0C, 0x18, 0x08, 0x2E, 0x4A, 0x37, 0x29, 0x03, 0x23,
	0x31, 0x3E, 0x3A, 0x38, 0x02, 0x11, 0x04, 0x5F, 0x72, 0x1D, 0x0C, 0x06,
	0x1F, 0x20, 0x19, 0x2F, 0x0F, 0x3E, 0x27, 0x16, 0x0E, 0x3C, 0x26, 0x34,
	0x28, 0x04, 0x21, 0x1F, 0x21, 0x22, 0x03, 0x2A, 0x59, 0x03, 0x22, 0x4A,
	0x5A, 0x26, 0x03, 0x20, 0x2A, 0x0B, 0x3F, 0x0B, 0x28, 0x2B, 0x02, 0x1E,
	0x2F, 0x39, 0x50, 0x01, 0x5C, 0x0B, 0x25, 0x36, 0x34, 0x33, 0x76, 0x2A,
	0x11, 0x25, 0x1F, 0x38, 0x06, 0x0B, 0x26, 0x0F, 0x7A, 0x38, 0x16, 0x0F,
	0x11, 0x6D, 0x19, 0x30, 0x1E, 0x2D, 0x0C, 0x3F, 0x03, 0x56, 0x32, 0x23,
	0x59, 0x58, 0x2D, 0x58, 0x07, 0x04, 0x11, 0x02, 0x22, 0x36, 0x54, 0x03,
	0x5B, 0x13, 0x0A, 0x59, 0x57, 0x09, 0x53, 0x35, 0x54, 0x15, 0x5D, 0x52,
	0x07, 0x3E, 0x25, 0x34, 0x09, 0x14, 0x2D, 0x20, 0x5E, 0x23, 0x03, 0x09,
	0x23, 0x56, 0x40, 0x0F, 0x58, 0x55, 0x26, 0x01, 0x18, 0x55, 0x10, 0x08,
	0x2D, 0x35, 0x1E, 0x03, 0x1F, 0x0C, 0x30, 0x43, 0x17, 0x27, 0x1C, 0x0D,
	0x18, 0x17, 0x3B, 0x2A, 0x25, 0x19, 0x15, 0x2D, 0x25, 0x24, 0x28, 0x39,
	0x1F, 0x06, 0x10, 0x23, 0x06, 0x3D, 0x3A, 0x2E, 0x14, 0x16, 0x18, 0x08,
	0x35, 0x34, 0x31, 0x27, 0x26, 0x17, 0x24, 0x2B, 0x0B, 0x59, 0x76, 0x09,
	0x07, 0x18, 0x33, 0x06, 0x0F, 0x00, 0x0B, 0x05, 0x70, 0x36, 0x24, 0x0F,
	0x11, 0x01, 0x3D, 0x59, 0x37, 0x1F, 0x21, 0x1F, 0x2F, 0x2C, 0x24, 0x12,
	0x22, 0x05, 0x5E, 0x5C, 0x28, 0x5B, 0x25, 0x0D, 0x08, 0x16, 0x24, 0x04,
	0x5C, 0x40, 0x16, 0x35, 0x0C, 0x45, 0x5B, 0x0E, 0x0A, 0x23, 0x14, 0x13,
	0x13, 0x5F, 0x08, 0x20, 0x05, 0x35, 0x0D, 0x20, 0x28, 0x20, 0x15, 0x3C,
	0x12, 0x29, 0x39, 0x33, 0x28, 0x11, 0x36, 0x08, 0x75, 0x18, 0x18, 0x07,
	0x5E, 0x03, 0x15, 0x23, 0x5B, 0x06, 0x12, 0x23, 0x26, 0x5A, 0x3E, 0x35,
	0x38, 0x26, 0x5A, 0x2E, 0x2D, 0x00, 0x02, 0x20, 0x2D, 0x16, 0x39, 0x04,
	0x03, 0x2E, 0x0D, 0x27, 0x11, 0x14, 0x26, 0x08, 0x38, 0x2F, 0x1D, 0x31,
	0x38, 0x47, 0x2F, 0x24, 0x5D, 0x0A, 0x26, 0x29, 0x3A, 0x5B, 0x23, 0x0B,
	0x1B, 0x5D, 0x5A, 0x0A, 0x23, 0x31, 0x19, 0x5D, 0x21, 0x20, 0x08, 0x3E,
	0x1D, 0x09, 0x04, 0x0E, 0x34, 0x2F, 0x33, 0x55, 0x14, 0x2B, 0x25, 0x1B,
	0x59, 0x58, 0x39, 0x1C, 0x03, 0x25, 0x58, 0x3A, 0x12, 0x6D, 0x1B, 0x22,
	0x14, 0x22, 0x0F, 0x36, 0x31, 0x27, 0x01, 0x2C, 0x03, 0x4E, 0x5A, 0x28,
	0x0A, 0x5B, 0x51, 0x0A, 0x53, 0x24, 0x24, 0x58, 0x1B, 0x3D, 0x04, 0x54,
	0x2F, 0x27, 0x52, 0x11, 0x2F, 0x0F, 0x59, 0x3D, 0x0E, 0x19, 0x53, 0x0D,
	0x18, 0x30, 0x58, 0x0B, 0x3F, 0x01, 0x23, 0x27, 0x18, 0x03, 0x20, 0x05,
	0x07, 0x28, 0x0B, 0x08, 0x20, 0x5D, 0x07, 0x17, 0x0F, 0x71, 0x05, 0x50,
	0x5A, 0x2F, 0x70, 0x59, 0x20, 0x0B, 0x1C, 0x00, 0x0E, 0x16, 0x3F, 0x05,
	0x0E, 0x43, 0x00, 0x29, 0x08, 0x24, 0x20, 0x15, 0x37, 0x04, 0x23, 0x26,
	0x57, 0x1B, 0x0F, 0x0C, 0x04, 0x29, 0x34, 0x3B, 0x35, 0x3D, 0x28, 0x03,
	0x11, 0x36, 0x29, 0x2E, 0x5E, 0x1B, 0x1A, 0x38, 0x12, 0x3D, 0x24, 0x69,
	0x09, 0x08, 0x59, 0x1A, 0x77, 0x0E, 0x52, 0x00, 0x5F, 0x32, 0x3F, 0x55,
	0x45, 0x28, 0x2F, 0x18, 0x0C, 0x3B, 0x1D, 0x37, 0x1E, 0x18, 0x03, 0x0C,
	0x11, 0x02, 0x32, 0x08, 0x38, 0x3B, 0x1E, 0x36, 0x0D, 0x3E, 0x15, 0x1A,
	0x2C, 0x3D, 0x52, 0x73, 0x5C, 0x0B, 0x0D, 0x5D, 0x6D, 0x20, 0x2D, 0x3D,
	0x32, 0x12, 0x3F, 0x0B, 0x1F, 0x01, 0x33, 0x23, 0x0D, 0x29, 0x0A, 0x73,
	0x06, 0x0B, 0x16, 0x39, 0x08, 0x55, 0x50, 0x09, 0x33, 0x14, 0x35, 0x26,
	0x28, 0x1E, 0x09, 0x36, 0x24, 0x26, 0x53, 0x0C, 0x55, 0x2F, 0x14, 0x18,
	0x75, 0x2E, 0x0F, 0x41, 0x52, 0x11, 0x06, 0x06, 0x05, 0x59, 0x75, 0x0F,
	0x22, 0x26, 0x1F, 0x26, 0x25, 0x05, 0x08, 0x28, 0x75, 0x03, 0x16, 0x39,
	0x1F, 0x28, 0x5D, 0x50, 0x1D, 0x5B, 0x32, 0x1F, 0x05, 0x3D, 0x5F, 0x72,
	0x29, 0x58, 0x17, 0x22, 0x7A, 0x38, 0x2C, 0x25, 0x0F, 0x27, 0x19, 0x2E,
	0x0A, 0x05, 0x34, 0x15, 0x00, 0x5C, 0x28, 0x1A, 0x06, 0x59, 0x34, 0x0D,
	0x7B, 0x55, 0x25, 0x06, 0x0D, 0x28, 0x2F, 0x27, 0x18, 0x59, 0x01, 0x5E,
	0x0F, 0x1B, 0x1D, 0x00, 0x1C, 0x59, 0x17, 0x06, 0x31, 0x5E, 0x0F, 0x17,
	0x5A, 0x25, 0x27, 0x54, 0x5D, 0x3B, 0x29, 0x21, 0x19, 0x1D, 0x1D, 0x16,
	0x22, 0x24, 0x19, 0x09, 0x31, 0x18, 0x27, 0x5B, 0x3E, 0x14, 0x36, 0x59,
	0x27, 0x09, 0x11, 0x22, 0x07, 0x2B, 0x05, 0x31, 0x35, 0x07, 0x19, 0x2C,
	0x29, 0x04, 0x19, 0x00, 0x5F, 0x23, 0x0F, 0x04, 0x26, 0x1D, 0x23, 0x04,
	0x14, 0x3D, 0x52, 0x23, 0x47, 0x28, 0x03, 0x3A, 0x17, 0x55, 0x33, 0x20,
	0x44, 0x27, 0x1C, 0x50, 0x39, 0x1D, 0x7B, 0x04, 0x2C, 0x22, 0x1C, 0x0A,
	0x5F, 0x25, 0x2D, 0x01, 0x11, 0x1B, 0x26, 0x57, 0x5E, 0x16, 0x3A, 0x06,
	0x14, 0x01, 0x2D, 0x21, 0x06, 0x28, 0x18, 0x18, 0x47, 0x23, 0x5E, 0x5B,
	0x2A, 0x0A, 0x38, 0x3F, 0x21, 0x2F, 0x09, 0x35, 0x36, 0x3F, 0x3B, 0x0F,
	0x17, 0x37, 0x59, 0x0A, 0x18, 0x51, 0x2F, 0x13, 0x0F, 0x3A, 0x53, 0x21,
	0x29, 0x21, 0x54, 0x11, 0x16, 0x0C, 0x26, 0x3B, 0x0E, 0x0A, 0x23, 0x12,
	0x0E, 0x52, 0x16, 0x29, 0x38, 0x5B, 0x20, 0x09, 0x02, 0x20, 0x0D, 0x53,
	0x45, 0x59, 0x27, 0x2A, 0x56, 0x17, 0x3C, 0x7B, 0x59, 0x0F, 0x1D, 0x2F,
	0x2B, 0x3A, 0x0C, 0x00, 0x28, 0x20, 0x06, 0x02, 0x2A, 0x3D, 0x25, 0x35,
	0x31, 0x56, 0x3C, 0x2B, 0x5E, 0x18, 0x5B, 0x0A, 0x28, 0x03, 0x17, 0x2D,
	0x0F, 0x16, 0x18, 0x27, 0x45, 0x1B, 0x76, 0x06, 0x08, 0x2F, 0x38, 0x74,
	0x22, 0x05, 0x2C, 0x38, 0x06, 0x01, 0x0F, 0x5F, 0x12, 0x75, 0x29, 0x08,
	0x41, 0x39, 0x77, 0x3E, 0x0B, 0x57, 0x03, 0x74, 0x55, 0x26, 0x1D, 0x32,
	0x1A, 0x3F, 0x36, 0x1B, 0x5C, 0x70, 0x54, 0x34, 0x34, 0x23, 0x16, 0x0F,
	0x0A, 0x37, 0x13, 0x2A, 0x14, 0x15, 0x1B, 0x40, 0x18, 0x18, 0x32, 0x57,
	0x2F, 0x2A, 0x20, 0x19, 0x03, 0x5C, 0x2A, 0x58, 0x19, 0x0C, 0x05, 0x01,
	0x1E, 0x54, 0x58, 0x24, 0x69, 0x14, 0x31, 0x56, 0x5F, 0x2B, 0x16, 0x2F,
	0x0D, 0x07, 0x29, 0x15, 0x29, 0x3A, 0x52, 0x35, 0x05, 0x4E, 0x0D, 0x25,
	0x29, 0x3C, 0x54, 0x19, 0x0A, 0x06, 0x43, 0x30, 0x3B, 0x1F, 0x0C, 0x2F,
	0x2B, 0x24, 0x28, 0x00, 0x2B, 0x1B, 0x5C, 0x0A, 0x26, 0x35, 0x53, 0x25,
	0x1A, 0x32, 0x26, 0x3B, 0x5B, 0x02, 0x04, 0x15, 0x17, 0x3B, 0x27, 0x08,
	0x1D, 0x52, 0x58, 0x29, 0x3B, 0x24, 0x36, 0x19, 0x00, 0x30, 0x22, 0x2E,
	0x1E, 0x06, 0x73, 0x09, 0x35, 0x16, 0x26, 0x24, 0x55, 0x0E, 0x1D, 0x12,
	0x37, 0x1E, 0x52, 0x03, 0x21, 0x04, 0x24, 0x0B, 0x24, 0x12, 0x7A, 0x1B,
	0x00, 0x04, 0x1C, 0x35, 0x1F, 0x37, 0x3C, 0x21, 0x24, 0x3A, 0x07, 0x29,
	0x1C, 0x00, 0x1D, 0x34, 0x34, 0x3E, 0x73, 0x03, 0x4E, 0x01, 0x5A, 0x69,
	0x02, 0x51, 0x04, 0x5C, 0x03, 0x35, 0x58, 0x03, 0x13, 0x06, 0x5F, 0x23,
	0x57, 0x1E, 0x2B, 0x24, 0x17, 0x05, 0x28, 0x0D, 0x20, 0x07, 0x5A, 0x2D,
	0x10, 0x21, 0x56, 0x59, 0x33, 0x76, 0x04, 0x25, 0x14, 0x1D, 0x13, 0x34,
	0x36, 0x29, 0x2F, 0x06, 0x14, 0x2D, 0x45, 0x03, 0x36, 0x14, 0x02, 0x59,
	0x5F, 0x24, 0x55, 0x18, 0x3E, 0x3B, 0x6D, 0x43, 0x56, 0x39, 0x44, 0x77,
	0x0A, 0x18, 0x3A, 0x22, 0x76, 0x3E, 0x52, 0x56, 0x11, 0x0D, 0x39, 0x12,
	0x5B, 0x27, 0x2A, 0x5B, 0x54, 0x3A, 0x29, 0x73, 0x5D, 0x02, 0x01, 0x39,
	0x29, 0x00, 0x12, 0x39, 0x38, 0x21, 0x15, 0x38, 0x1E, 0x21, 0x04, 0x0F,
	0x56, 0x07, 0x2E, 0x05, 0x54, 0x32, 0x2B, 0x3E, 0x2F, 0x01, 0x19, 0x56,
	0x12, 0x21, 0x5C, 0x38, 0x14, 0x2A, 0x0D, 0x58, 0x29, 0x56, 0x52, 0x1B,
	0x5A, 0x03, 0x1A, 0x11, 0x21, 0x2A, 0x11, 0x14, 0x5E, 0x20, 0x04, 0x11,
	0x5D, 0x38, 0x2A, 0x1E, 0x38, 0x06, 0x20, 0x12, 0x04, 0x04, 0x23, 0x52,
	0x24, 0x24, 0x2E, 0x27, 0x2A, 0x32, 0x5A, 0x3B, 0x2B, 0x5D, 0x05, 0x2D,
	0x24, 0x5A, 0x1F, 0x73, 0x24, 0x27, 0x59, 0x1F, 0x1A, 0x35, 0x22, 0x07,
	0x3E, 0x28, 0x47, 0x2F, 0x2D, 0x20, 0x2B, 0x02, 0x16, 0x05, 0x1F, 0x38,
	0x01, 0x2B, 0x28, 0x44, 0x01, 0x3C, 0x0E, 0x04, 0x3F, 0x75, 0x43, 0x02,
	0x5E, 0x1E, 0x07, 0x2F, 0x14, 0x25, 0x0C, 0x6D, 0x5C, 0x26, 0x3D, 0x09,
	0x13, 0x5F, 0x19, 0x56, 0x13, 0x06, 0x5B, 0x18, 0x25, 0x1D, 0x14, 0x3E,
	0x14, 0x59, 0x5B, 0x0A, 0x26, 0x2D, 0x0A, 0x29, 0x31, 0x15, 0x12, 0x38,
	0x0D, 0x33, 0x09, 0x2D, 0x3E, 0x23, 0x73, 0x20, 0x27, 0x0C, 0x5C, 0x27,
	0x14, 0x05, 0x1C, 0x2D, 0x21, 0x2A, 0x06, 0x02, 0x0F, 0x24, 0x55, 0x12,
	0x1A, 0x06, 0x76, 0x23, 0x05, 0x2A, 0x5E, 0x12, 0x5F, 0x57, 0x1A, 0x01,
	0x31, 0x34, 0x39, 0x1F, 0x0F, 0x2C, 0x26, 0x19, 0x58, 0x3E, 0x32, 0x1B,
	0x26, 0x5F, 0x59, 0x26, 0x54, 0x33, 0x5A, 0x1E, 0x18, 0x1F, 0x56, 0x1C,
	0x27, 0x2C, 0x0D, 0x53, 0x19, 0x5C, 0x0D, 0x39, 0x29, 0x36, 0x5E, 0x6D,
	0x07, 0x26, 0x0F, 0x38, 0x2E, 0x5C, 0x14, 0x14, 0x0D, 0x2F, 0x5D, 0x2E,
	0x5D, 0x20, 0x38, 0x1A, 0x0F, 0x23, 0x26, 0x15, 0x54, 0x53, 0x26, 0x1F,
	0x71, 0x22, 0x53, 0x41, 0x33, 0x7A, 0x43, 0x56, 0x34, 0x1D, 0x6D, 0x43,
	0x17, 0x34, 0x5D, 0x34, 0x16, 0x02, 0x3A, 0x5A, 0x75, 0x28, 0x2C, 0x00,
	0x1D, 0x0A, 0x38, 0x57, 0x21, 0x31, 0x0A, 0x5D, 0x4E, 0x26, 0x5A, 0x70,
	0x23, 0x31, 0x26, 0x59, 0x08, 0x5B, 0x35, 0x5F, 0x0D, 0x01, 0x06, 0x28,
	0x0C, 0x02, 0x71, 0x22, 0x30, 0x1F, 0x5F, 0x15, 0x5F, 0x24, 0x2F, 0x38,
	0x38, 0x43, 0x51, 0x25, 0x28, 0x27, 0x14, 0x14, 0x23, 0x11, 0x05, 0x27,
	0x28, 0x26, 0x3B, 0x26, 0x54, 0x4A, 0x09, 0x07, 0x10, 0x5A, 0x04, 0x24,
	0x40, 0x73, 0x01, 0x34, 0x06, 0x26, 0x21, 0x35, 0x35, 0x5D, 0x1F, 0x37,
	0x28, 0x50, 0x2A, 0x39, 0x3B, 0x02, 0x05, 0x2F, 0x3F, 0x29, 0x58, 0x28,
	0x5D, 0x5A, 0x31, 0x2D, 0x10, 0x0A, 0x32, 0x7B, 0x35, 0x05, 0x07, 0x52,
	0x10, 0x5C, 0x57, 0x5F, 0x25, 0x21, 0x54, 0x09, 0x59, 0x2A, 0x0E, 0x24,
	0x35, 0x1F, 0x3B, 0x7A, 0x5D, 0x0D, 0x1C, 0x3B, 0x2D, 0x08, 0x38, 0x41,
	0x03, 0x3A, 0x16, 0x27, 0x45, 0x3B, 0x28, 0x16, 0x54, 0x2D, 0x5A, 0x3A,
	0x28, 0x59, 0x2D, 0x3C, 0x2F, 0x5D, 0x0B, 0x22, 0x2A, 0x6D, 0x0F, 0x30,
	0x1A, 0x5C, 0x35, 0x24, 0x53, 0x45, 0x5E, 0x05, 0x3D, 0x0F, 0x1C, 0x00,
	0x20, 0x24, 0x03, 0x34, 0x53, 0x0F, 0x5F, 0x51, 0x34, 0x05, 0x2F, 0x09,
	0x2D, 0x0A, 0x5B, 0x0F, 0x1A, 0x32, 0x37, 0x0D, 0x05, 0x38, 0x50, 0x45,
	0x40, 0x11, 0x09, 0x05, 0x2A, 0x11, 0x7B, 0x02, 0x2F, 0x1E, 0x5B, 0x12,
	0x08, 0x19, 0x5A, 0x22, 0x06, 0x2B, 0x18, 0x04, 0x00, 0x0A, 0x2E, 0x39,
	0x36, 0x07, 0x27, 0x03, 0x0E, 0x2C, 0x0D, 0x21, 0x36, 0x58, 0x28, 0x03,
	0x2C, 0x21, 0x1B, 0x41, 0x27, 0x31, 0x3C, 0x25, 0x21, 0x26, 0x75, 0x14,
	0x0E, 0x02, 0x20, 0x1B, 0x27, 0x29, 0x1C, 0x11, 0x38, 0x02, 0x0A, 0x0B,
	0x32, 0x69, 0x23, 0x0F, 0x24, 0x00, 0x30, 0x09, 0x09, 0x34, 0x2E, 0x0E,
	0x2A, 0x05, 0x57, 0x07, 0x7A, 0x18, 0x53, 0x1B, 0x0F, 0x09, 0x3B, 0x1B,
	0x21, 0x23, 0x25, 0x08, 0x33, 0x0D, 0x0F, 0x34, 0x2D, 0x59, 0x3C, 0x1F,
	0x25, 0x5C, 0x10, 0x2F, 0x11, 0x08, 0x5B, 0x0F, 0x21, 0x5C, 0x69, 0x1A,
	0x2F, 0x3B, 0x1D, 0x07, 0x09, 0x58, 0x59, 0x1B, 0x06, 0x24, 0x07, 0x3B,
	0x27, 0x12, 0x34, 0x0B, 0x45, 0x3C, 0x2D, 0x00, 0x53, 0x3D, 0x0A, 0x24,
	0x0B, 0x56, 0x0D, 0x08, 0x33, 0x0B, 0x2C, 0x05, 0x1C, 0x12, 0x58, 0x39,
	0x01, 0x52, 0x69, 0x22, 0x22, 0x38, 0x09, 0x28, 0x43, 0x12, 0x3C, 0x1E,
	0x03, 0x3C, 0x26, 0x1A, 0x04, 0x05, 0x1F, 0x26, 0x58, 0x20, 0x18, 0x1E,
	0x37, 0x5C, 0x3C, 0x2B, 0x24, 0x34, 0x21, 0x0C, 0x08, 0x18, 0x23, 0x0B,
	0x5B, 0x10, 0x1D, 0x1B, 0x14, 0x33, 0x08, 0x35, 0x59, 0x28, 0x13, 0x00,
	0x08, 0x14, 0x0A, 0x2A, 0x06, 0x54, 0x56, 0x3F, 0x18, 0x77, 0x2F, 0x4A,
	0x2A, 0x05, 0x2C, 0x06, 0x0B, 0x23, 0x01, 0x7B, 0x04, 0x58, 0x1A, 0x5B,
	0x1A, 0x29, 0x26, 0x29, 0x02, 0x34, 0x0F, 0x07, 0x37, 0x02, 0x31, 0x00,
	0x53, 0x04, 0x00, 0x3A, 0x2D, 0x12, 0x01, 0x13, 0x0C, 0x1B, 0x24, 0x02,
	0x02, 0x20, 0x38, 0x06, 0x14, 0x21, 0x27, 0x3B, 0x19, 0x09, 0x2D, 0x04,
	0x5B, 0x53, 0x05, 0x3B, 0x04, 0x21, 0x07, 0x5E, 0x02, 0x23, 0x39, 0x2C,
	0x26, 0x04, 0x77, 0x24, 0x4E, 0x09, 0x2E, 0x15, 0x19, 0x23, 0x41, 0x44,
	0x36, 0x23, 0x05, 0x08, 0x0D, 0x01, 0x09, 0x23, 0x04, 0x1B, 0x28, 0x24,
	0x39, 0x5C, 0x00, 0x15, 0x2D, 0x34, 0x04, 0x12, 0x23, 0x2D, 0x25, 0x27,
	0x3B, 0x05, 0x5F, 0x2E, 0x3A, 0x00, 0x7B, 0x07, 0x17, 0x00, 0x0D, 0x11,
	0x0A, 0x29, 0x20, 0x04, 0x7A, 0x26, 0x56, 0x1E, 0x1B, 0x71, 0x2B, 0x4A,
	0x57, 0x5B, 0x72, 0x3C, 0x1B, 0x5D, 0x0F, 0x12, 0x3D, 0x52, 0x07, 0x40,
	0x03, 0x55, 0x57, 0x2D, 0x40, 0x26, 0x59, 0x1B, 0x21, 0x05, 0x35, 0x3C,
	0x09, 0x2D, 0x05, 0x06, 0x38, 0x07, 0x17, 0x06, 0x36, 0x16, 0x17, 0x2D,
	0x09, 0x70, 0x36, 0x4E, 0x2D, 0x03, 0x09, 0x5F, 0x08, 0x2F, 0x29, 0x2F,
	0x26, 0x14, 0x41, 0x3B, 0x2F, 0x1F, 0x23, 0x18, 0x31, 0x03, 0x1E, 0x50,
	0x5F, 0x1F, 0x75, 0x5E, 0x2C, 0x57, 0x33, 0x38, 0x5C, 0x0A, 0x34, 0x32,
	0x2A, 0x22, 0x0E, 0x5D, 0x5B, 0x16, 0x38, 0x55, 0x19, 0x08, 0x71, 0x1F,
	0x0D, 0x20, 0x25, 0x2D, 0x20, 0x20, 0x1C, 0x26, 0x1A, 0x29, 0x56, 0x29,
	0x5C, 0x05, 0x54, 0x19, 0x03, 0x58, 0x6D, 0x24, 0x1B, 0x08, 0x2F, 0x3B,
	0x0F, 0x03, 0x17, 0x53, 0x1B, 0x3E, 0x26, 0x5E, 0x58, 0x0C, 0x24, 0x07,
	0x00, 0x5B, 0x09, 0x24, 0x0F, 0x5B, 0x44, 0x0D, 0x07, 0x12, 0x0B, 0x07,
	0x25, 0x20, 0x11, 0x01, 0x1E, 0x16, 0x2A, 0x33, 0x0D, 0x2D, 0x7B, 0x26,
	0x03, 0x23, 0x38, 0x23, 0x20, 0x12, 0x1F, 0x0E, 0x27, 0x06, 0x10, 0x0B,
	0x5C, 0x2E, 0x29, 0x11, 0x1E, 0x2A, 0x2C, 0x1B, 0x35, 0x07, 0x20, 0x35,
	0x06, 0x25, 0x0C, 0x01, 0x7B, 0x59, 0x2C, 0x28, 0x0F, 0x74, 0x5A, 0x04,
	0x37, 0x59, 0x21, 0x28, 0x18, 0x27, 0x52, 0x33, 0x5E, 0x32, 0x14, 0x26,
	0x69, 0x03, 0x24, 0x1D, 0x13, 0x24, 0x18, 0x35, 0x3C, 0x22, 0x1A, 0x1D,
	0x55, 0x29, 0x59, 0x23, 0x1F, 0x50, 0x3D, 0x26, 0x06, 0x15, 0x50, 0x23,
	0x18, 0x1B, 0x15, 0x24, 0x1E, 0x02, 0x6D, 0x29, 0x52, 0x01, 0x32, 0x18,
	0x38, 0x33, 0x0B, 0x29, 0x06, 0x02, 0x22, 0x24, 0x5E, 0x0F, 0x5C, 0x03,
	0x08, 0x29, 0x0A, 0x5A, 0x03, 0x59, 0x12, 0x0C, 0x39, 0x25, 0x0C, 0x18,
	0x70, 0x2B, 0x58, 0x02, 0x53, 0x35, 0x39, 0x05, 0x1C, 0x1B, 0x07, 0x5A,
	0x2F, 0x58, 0x1A, 0x06, 0x0B, 0x22, 0x14, 0x5E, 0x13, 0x3A, 0x23, 0x17,
	0x04, 0x0B, 0x2B, 0x59, 0x5C, 0x0C, 0x20, 0x2E, 0x0A, 0x5E, 0x0A, 0x28,
	0x16, 0x0B, 0x05, 0x5B, 0x01, 0x2D, 0x14, 0x17, 0x5F, 0x14, 0x01, 0x00,
	0x1A, 0x2D, 0x01, 0x28, 0x38, 0x3D, 0x25, 0x16, 0x2E, 0x2F, 0x0A, 0x13,
	0x10, 0x05, 0x4A, 0x25, 0x0A, 0x26, 0x35, 0x2C, 0x5A, 0x1F, 0x34, 0x02,
	0x2A, 0x08, 0x11, 0x76, 0x2B, 0x02, 0x3C, 0x1B, 0x69, 0x58, 0x25, 0x07,
	0x40, 0x27, 0x0F, 0x06, 0x0C, 0x3C, 0x24, 0x14, 0x22, 0x19, 0x3B, 0x20,
	0x00, 0x19, 0x3A, 0x07, 0x1B, 0x1E, 0x2F, 0x01, 0x40, 0x13, 0x58, 0x03,
	0x2B, 0x07, 0x3A, 0x58, 0x31, 0x36, 0x21, 0x76, 0x1B, 0x20, 0x01, 0x03,
	0x3B, 0x54, 0x51, 0x1E, 0x04, 0x2F, 0x39, 0x4A, 0x34, 0x03, 0x20, 0x3C,
	0x06, 0x21, 0x5F, 0x0B, 0x27, 0x20, 0x00, 0x53, 0x69, 0x2D, 0x19, 0x1D,
	0x1B, 0x09, 0x02, 0x0E, 0x3B, 0x3F, 0x30, 0x43, 0x04, 0x38, 0x3A, 0x26,
	0x0B, 0x52, 0x08, 0x33, 0x09, 0x3F, 0x2F, 0x06, 0x5C, 0x28, 0x55, 0x32,
	0x07, 0x32, 0x35, 0x3B, 0x12, 0x39, 0x39, 0x73, 0x2F, 0x15, 0x41, 0x24,
	0x74, 0x5A, 0x17, 0x0A, 0x25, 0x3A, 0x2D, 0x31, 0x27, 0x52, 0x21, 0x23,
	0x39, 0x28, 0x00, 0x0F, 0x00, 0x15, 0x06, 0x26, 0x12, 0x05, 0x15, 0x18,
	0x3B, 0x26, 0x02, 0x58, 0x1B, 0x52, 0x1A, 0x38, 0x17, 0x5A, 0x2C, 0x35,
	0x47, 0x22, 0x14, 0x59, 0x6D, 0x2E, 0x16, 0x20, 0x2A, 0x73, 0x0E, 0x54,
	0x24, 0x1F, 0x03, 0x5A, 0x50, 0x2C, 0x53, 0x1A, 0x35, 0x2B, 0x0D, 0x58,
	0x32, 0x1B, 0x32, 0x03, 0x0A, 0x24, 0x09, 0x12, 0x3D, 0x3E, 0x33, 0x14,
	0x36, 0x38, 0x22, 0x05, 0x5D, 0x0B, 0x17, 0x27, 0x12, 0x1A, 0x04, 0x56,
	0x3F, 0x13, 0x22, 0x54, 0x14, 0x06, 0x20, 0x36, 0x54, 0x2B, 0x02, 0x0C,
	0x1B, 0x23, 0x34, 0x26, 0x1A, 0x5E, 0x17, 0x01, 0x31, 0x72, 0x02, 0x2E,
	0x0B, 0x3C, 0x17, 0x0B, 0x30, 0x07, 0x5C, 0x2C, 0x05, 0x55, 0x26, 0x00,
	0x2C, 0x2A, 0x59, 0x22, 0x2F, 0x3A, 0x0D, 0x52, 0x1F, 0x07, 0x35, 0x1C,
	0x04, 0x1F, 0x40, 0x12, 0x1E, 0x0A, 0x38, 0x5F, 0x20, 0x39, 0x28, 0x41,
	0x3C, 0x7B, 0x29, 0x39, 0x3D, 0x12, 0x69, 0x5C, 0x22, 0x1C, 0x2A, 0x37,
	0x35, 0x16, 0x0F, 0x38, 0x7B, 0x55, 0x36, 0x16, 0x3B, 0x34, 0x2E, 0x00,
	0x39, 0x44, 0x10, 0x5B, 0x0E, 0x27, 0x1E, 0x20, 0x27, 0x31, 0x37, 0x26,
	0x17, 0x29, 0x35, 0x16, 0x25, 0x0F, 0x3A, 0x06, 0x04, 0x5F, 0x18, 0x20,
	0x08, 0x2A, 0x0E, 0x27, 0x27, 0x15, 0x1F, 0x27, 0x23, 0x15, 0x31, 0x3B,
	0x1A, 0x17, 0x3B, 0x2C, 0x29, 0x1B, 0x23, 0x38, 0x06, 0x2F, 0x25, 0x10,
	0x2E, 0x10, 0x0F, 0x1C, 0x25, 0x36, 0x17, 0x09, 0x11, 0x1A, 0x2A, 0x53,
	0x14, 0x28, 0x2A, 0x1B, 0x50, 0x25, 0x20, 0x21, 0x54, 0x53, 0x1D, 0x0A,
	0x06, 0x0E, 0x02, 0x08, 0x31, 0x05, 0x1A, 0x52, 0x07, 0x02, 0x32, 0x34,
	0x33, 0x1B, 0x0D, 0x2F, 0x0A, 0x30, 0x24, 0x0C, 0x04, 0x01, 0x23, 0x04,
	0x07, 0x27, 0x38, 0x2C, 0x1C, 0x52, 0x0D, 0x05, 0x26, 0x21, 0x3B, 0x1B,
	0x29, 0x0B, 0x09, 0x20, 0x2C, 0x36, 0x38, 0x07, 0x58, 0x01, 0x34, 0x2D,
	0x16, 0x59, 0x3B, 0x08, 0x34, 0x45, 0x03, 0x38, 0x18, 0x25, 0x2D, 0x0E,
	0x05, 0x1B, 0x23, 0x1C, 0x2A, 0x7A, 0x43, 0x0B, 0x41, 0x0E, 0x14, 0x03,
	0x05, 0x5E, 0x5B, 0x28, 0x1A, 0x02, 0x2D, 0x39, 0x32, 0x04, 0x08, 0x26,
	0x3F, 0x09, 0x3C, 0x38, 0x04, 0x58, 0x74, 0x2D, 0x2C, 0x0B, 0x3D, 0x32,
	0x2B, 0x12, 0x34, 0x08, 0x18, 0x35, 0x06, 0x57, 0x23, 0x3A, 0x01, 0x1B,
	0x04, 0x1A, 0x0E, 0x54, 0x13, 0x24, 0x05, 0x15, 0x21, 0x0E, 0x1D, 0x59,
	0x2F, 0x29, 0x57, 0x25, 0x07, 0x2A, 0x0E, 0x23, 0x57, 0x38, 0x27, 0x05,
	0x51, 0x1D, 0x03, 0x07, 0x3F, 0x53, 0x29, 0x20, 0x76, 0x28, 0x26, 0x3F,
	0x5D, 0x77, 0x3B, 0x36, 0x20, 0x1F, 0x01, 0x05, 0x59, 0x37, 0x2C, 0x18,
	0x38, 0x16, 0x41, 0x01, 0x00, 0x3C, 0x05, 0x21, 0x39, 0x2C, 0x28, 0x54,
	0x59, 0x3A, 0x2A, 0x23, 0x26, 0x3D, 0x5B, 0x01, 0x1E, 0x35, 0x19, 0x2D,
	0x74, 0x02, 0x4A, 0x3C, 0x2E, 0x1A, 0x59, 0x2C, 0x22, 0x08, 0x23, 0x5B,
	0x0A, 0x02, 0x18, 0x18, 0x2E, 0x38, 0x58, 0x29, 0x2A, 0x2A, 0x17, 0x2A,
	0x24, 0x24, 0x08, 0x30, 0x04, 0x1B, 0x2C, 0x5C, 0x0C, 0x20, 0x2C, 0x71,
	0x3D, 0x34, 0x24, 0x0E, 0x0D, 0x27, 0x04, 0x2F, 0x08, 0x32, 0x1C, 0x3B,
	0x00, 0x0D, 0x05, 0x3D, 0x02, 0x29, 0x2E, 0x76, 0x59, 0x53, 0x22, 0x20,
	0x70, 0x0F, 0x23, 0x17, 0x23, 0x2D, 0x27, 0x24, 0x0C, 0x1E, 0x05, 0x0F,
	0x3B, 0x23, 0x19, 0x77, 0x0B, 0x2E, 0x38, 0x26, 0x25, 0x03, 0x30, 0x04,
	0x33, 0x70, 0x1F, 0x54, 0x14, 0x3E, 0x15, 0x35, 0x0A, 0x56, 0x1D, 0x74,
	0x01, 0x30, 0x01, 0x21, 0x34, 0x58, 0x33, 0x14, 0x0F, 0x2E, 0x2E, 0x2E,
	0x3A, 0x53, 0x32, 0x3E, 0x3B, 0x06, 0x22, 0x14, 0x2B, 0x11, 0x0B, 0x23,
	0x0F, 0x5F, 0x4A, 0x07, 0x11, 0x04, 0x5F, 0x34, 0x01, 0x2F, 0x09, 0x24,
	0x3B, 0x0C, 0x5F, 0x14, 0x16, 0x17, 0x17, 0x2A, 0x0F, 0x1C, 0x04, 0x19,
	0x11, 0x04, 0x27, 0x36, 0x21, 0x38, 0x0D, 0x0F, 0x57, 0x0F, 0x23, 0x0F,
	0x5E, 0x32, 0x16, 0x11, 0x03, 0x0F, 0x14, 0x56, 0x27, 0x77, 0x16, 0x54,
	0x2B, 0x2C, 0x1A, 0x09, 0x16, 0x3A, 0x22, 0x1A, 0x1F, 0x12, 0x17, 0x28,
	0x21, 0x23, 0x3B, 0x01, 0x12, 0x31, 0x14, 0x0A, 0x03, 0x32, 0x36, 0x35,
	0x54, 0x05, 0x33, 0x2A, 0x16, 0x22, 0x29, 0x3E, 0x3B, 0x0E, 0x29, 0x23,
	0x19, 0x73, 0x00, 0x0C, 0x57, 0x58, 0x00, 0x01, 0x2D, 0x56, 0x1B, 0x72,
	0x5C, 0x3B, 0x27, 0x04, 0x3B, 0x5D, 0x0F, 0x03, 0x04, 0x23, 0x55, 0x51,
	0x05, 0x2E, 0x18, 0x5F, 0x16, 0x2F, 0x1C, 0x38, 0x22, 0x0B, 0x5C, 0x2D,
	0x37, 0x02, 0x12, 0x14, 0x19, 0x08, 0x28, 0x57, 0x25, 0x52, 0x75, 0x02,
	0x02, 0x0C, 0x2A, 0x73, 0x59, 0x17, 0x5A, 0x0E, 0x32, 0x23, 0x24, 0x0B,
	0x09, 0x18, 0x2B, 0x27, 0x28, 0x1E, 0x14, 0x3B, 0x2F, 0x36, 0x08, 0x0A,
	0x1A, 0x06, 0x1F, 0x02, 0x7A, 0x04, 0x19, 0x0B, 0x3D, 0x69, 0x1F, 0x59,
	0x07, 0x23, 0x11, 0x08, 0x15, 0x07, 0x3B, 0x69, 0x02, 0x09, 0x5B, 0x0C,
	0x0C, 0x58, 0x20, 0x17, 0x12, 0x0A, 0x29, 0x59, 0x18, 0x13, 0x0B, 0x16,
	0x59, 0x14, 0x22, 0x17, 0x1E, 0x34, 0x34, 0x00, 0x33, 0x38, 0x16, 0x3A,
	0x01, 0x10, 0x08, 0x16, 0x5B, 0x0D, 0x2F, 0x01, 0x51, 0x5D, 0x5C, 0x70,
	0x1D, 0x27, 0x21, 0x0F, 0x75, 0x01, 0x02, 0x3E, 0x40, 0x3A, 0x39, 0x10,
	0x2A, 0x2F, 0x29, 0x3A, 0x17, 0x3F, 0x0E, 0x74, 0x23, 0x20, 0x36, 0x22,
	0x3B, 0x06, 0x4A, 0x28, 0x12, 0x05, 0x1E, 0x37, 0x2F, 0x2E, 0x16, 0x05,
	0x35, 0x34, 0x5A, 0x10, 0x00, 0x0C, 0x1D, 0x2A, 0x17, 0x36, 0x3B, 0x18,
	0x2A, 0x09, 0x43, 0x27, 0x5E, 0x3E, 0x24, 0x1C, 0x22, 0x06, 0x05, 0x01,
	0x5F, 0x4E, 0x2B, 0x29, 0x21, 0x39, 0x22, 0x37, 0x2F, 0x7A, 0x14, 0x13,
	0x04, 0x0E, 0x72, 0x5F, 0x2C, 0x2A, 0x29, 0x74, 0x1E, 0x50, 0x2D, 0x07,
	0x3A, 0x5F, 0x16, 0x25, 0x33, 0x21, 0x29, 0x38, 0x0F, 0x06, 0x04, 0x20,
	0x27, 0x1C, 0x58, 0x38, 0x01, 0x18, 0x09, 0x1A, 0x0C, 0x26, 0x14, 0x5B,
	0x31, 0x36, 0x1B, 0x4E, 0x0D, 0x03, 0x13, 0x07, 0x2C, 0x26, 0x53, 0x00,
	0x2A, 0x28, 0x25, 0x05, 0x18, 0x1B, 0x54, 0x59, 0x1D, 0x2E, 0x3C, 0x31,
	0x00, 0x1F, 0x76, 0x1D, 0x0C, 0x02, 0x29, 0x04, 0x2B, 0x38, 0x37, 0x1E,
	0x24, 0x3C, 0x16, 0x3F, 0x13, 0x26, 0x1C, 0x57, 0x56, 0x29, 0x1B, 0x35,
	0x25, 0x28, 0x2F, 0x13, 0x2D, 0x09, 0x3E, 0x06, 0x0E, 0x5E, 0x2B, 0x02,
	0x5A, 0x2F, 0x23, 0x3B, 0x0A, 0x5E, 0x1B, 0x38, 0x05, 0x2D, 0x0C, 0x11,
	0x2D, 0x37, 0x5A, 0x33, 0x16, 0x5E, 0x37, 0x38, 0x5E, 0x2D, 0x3F, 0x03,
	0x5E, 0x3E, 0x0B, 0x34, 0x31, 0x1F, 0x5E, 0x2B, 0x0E, 0x37, 0x2C, 0x26,
	0x35, 0x00, 0x4E, 0x2B, 0x22, 0x7A, 0x3E, 0x18, 0x22, 0x1C, 0x3A, 0x0E,
	0x00, 0x2C, 0x0E, 0x26, 0x0F, 0x2E, 0x1A, 0x1B, 0x20, 0x3A, 0x58, 0x1B,
	0x31, 0x0A, 0x1A, 0x10, 0x3C, 0x09, 0x2E, 0x1E, 0x16, 0x0B, 0x02, 0x01,
	0x59, 0x11, 0x23, 0x13, 0x69, 0x23, 0x29, 0x25, 0x5F, 0x74, 0x0D, 0x19,
	0x0B, 0x22, 0x16, 0x23, 0x50, 0x45, 0x44, 0x18, 0x5B, 0x33, 0x07, 0x3B,
	0x07, 0x2A, 0x0A, 0x41, 0x52, 0x26, 0x01, 0x15, 0x56, 0x2D, 0x76, 0x0F,
	0x14, 0x3C, 0x0F, 0x08, 0x0A, 0x33, 0x3A, 0x0D, 0x16, 0x5C, 0x07, 0x14,
	0x5C, 0x7A, 0x38, 0x52, 0x1D, 0x0A, 0x21, 0x06, 0x56, 0x58, 0x3B, 0x3A,
	0x43, 0x04, 0x22, 0x04, 0x69, 0x16, 0x23, 0x56, 0x5E, 0x74, 0x20, 0x17,
	0x02, 0x40, 0x06, 0x5B, 0x0D, 0x03, 0x01, 0x7B, 0x0F, 0x4E, 0x29, 0x52,
	0x0D, 0x36, 0x13, 0x08, 0x2A, 0x7B, 0x43, 0x39, 0x3C, 0x1F, 0x7B, 0x3C,
	0x03, 0x37, 0x23, 0x71, 0x18, 0x57, 0x3E, 0x1D, 0x13, 0x34, 0x19, 0x41,
	0x26, 0x34, 0x1D, 0x4A, 0x26, 0x0F, 0x7B, 0x24, 0x33, 0x20, 0x44, 0x1A,
	0x58, 0x56, 0x1D, 0x1B, 0x69, 0x1A, 0x55, 0x57, 0x1D, 0x33, 0x1A, 0x33,
	0x41, 0x01, 0x75, 0x24, 0x58, 0x5F, 0x3C, 0x10, 0x55, 0x4E, 0x0C, 0x40,
	0x00, 0x3C, 0x16, 0x45, 0x5A, 0x3A, 0x22, 0x57, 0x0A, 0x06, 0x3B, 0x03,
	0x36, 0x08, 0x38, 0x37, 0x3D, 0x11, 0x1D, 0x5C, 0x69, 0x59, 0x22, 0x38,
	0x11, 0x09, 0x15, 0x30, 0x58, 0x31, 0x2E, 0x05, 0x53, 0x03, 0x26, 0x2F,
	0x09, 0x27, 0x21, 0x08, 0x10, 0x3D, 0x03, 0x0C, 0x23, 0x69, 0x59, 0x39,
	0x09, 0x24, 0x07, 0x2D, 0x25, 0x38, 0x31, 0x1A, 0x04, 0x34, 0x59, 0x1F,
	0x26, 0x1B, 0x28, 0x41, 0x0C, 0x0E, 0x35, 0x26, 0x1A, 0x5F, 0x33, 0x18,
	0x30, 0x1D, 0x2E, 0x10, 0x0E, 0x3B, 0x20, 0x5F, 0x09, 0x1B, 0x3B, 0x22,
	0x02, 0x08, 0x35, 0x53, 0x34, 0x5F, 0x17, 0x1E, 0x35, 0x5D, 0x00, 0x05,
	0x5B, 0x4E, 0x39, 0x40, 0x30, 0x29, 0x07, 0x03, 0x52, 0x69, 0x0A, 0x1B,
	0x26, 0x24, 0x73, 0x3B, 0x31, 0x5F, 0x2E, 0x12, 0x1F, 0x15, 0x3F, 0x5D,
	0x03, 0x16, 0x29, 0x17, 0x1E, 0x11, 0x20, 0x02, 0x3E, 0x26, 0x38, 0x0F,
	0x02, 0x3C, 0x44, 0x12, 0x08, 0x35, 0x2A, 0x1A, 0x08, 0x2F, 0x4A, 0x08,
	0x1F, 0x03, 0x24, 0x34, 0x21, 0x0D, 0x30, 0x03, 0x36, 0x2F, 0x19, 0x15,
	0x1F, 0x03, 0x57, 0x2E, 0x36, 0x54, 0x52, 0x29, 0x13, 0x0B, 0x1A, 0x24,
	0x14, 0x5B, 0x21, 0x39, 0x17, 0x0F, 0x00, 0x00, 0x26, 0x52, 0x01, 0x1B,
	0x7A, 0x2F, 0x38, 0x1A, 0x0E, 0x10, 0x21, 0x28, 0x05, 0x06, 0x70, 0x3C,
	0x00, 0x14, 0x2E, 0x03, 0x04, 0x59, 0x3A, 0x20, 0x3B, 0x00, 0x25, 0x05,
	0x44, 0x0E, 0x05, 0x32, 0x04, 0x29, 0x04, 0x5A, 0x28, 0x2A, 0x39, 0x0A,
	0x0B, 0x00, 0x1E, 0x13, 0x31, 0x00, 0x06, 0x2F, 0x26, 0x2B, 0x5F, 0x14,
	0x22, 0x05, 0x29, 0x0A, 0x2C, 0x0A, 0x1D, 0x29, 0x02, 0x4E, 0x29, 0x3C,
	0x15, 0x02, 0x00, 0x0F, 0x04, 0x18, 0x2A, 0x58, 0x36, 0x5C, 0x1A, 0x0F,
	0x14, 0x38, 0x07, 0x72, 0x58, 0x00, 0x39, 0x2C, 0x3B, 0x55, 0x0F, 0x24,
	0x12, 0x1B, 0x1C, 0x34, 0x57, 0x2F, 0x04, 0x01, 0x2B, 0x1E, 0x12, 0x0A,
	0x59, 0x25, 0x5E, 0x1F, 0x0E, 0x3A, 0x04, 0x37, 0x0F, 0x16, 0x19, 0x26,
	0x08, 0x12, 0x32, 0x5E, 0x0B, 0x1B, 0x07, 0x32, 0x2A, 0x00, 0x3D, 0x0E,
	0x69, 0x3D, 0x39, 0x5D, 0x23, 0x2E, 0x25, 0x09, 0x45, 0x3B, 0x7A, 0x3A,
	0x24, 0x14, 0x1D, 0x76, 0x2F, 0x10, 0x18, 0x21, 0x17, 0x00, 0x11, 0x39,
	0x2F, 0x06, 0x1F, 0x0E, 0x3D, 0x2E, 0x31, 0x3C, 0x37, 0x3D, 0x1E, 0x04,
	0x24, 0x2F, 0x59, 0x13, 0x2E, 0x04, 0x36, 0x03, 0x53, 0x0B, 0x01, 0x11,
	0x3C, 0x24, 0x05, 0x2F, 0x0C, 0x59, 0x5C, 0x28, 0x25, 0x0D, 0x0B, 0x21,
	0x2E, 0x07, 0x11, 0x26, 0x3B, 0x6D, 0x1C, 0x0E, 0x3A, 0x3E, 0x38, 0x22,
	0x0A, 0x58, 0x2D, 0x33, 0x39, 0x02, 0x5A, 0x09, 0x00, 0x07, 0x39, 0x1A,
	0x04, 0x07, 0x38, 0x24, 0x34, 0x0F, 0x33, 0x25, 0x06, 0x5E, 0x28, 0x06,
	0x24, 0x3B, 0x18, 0x1E, 0x29, 0x0D, 0x0E, 0x16, 0x2F, 0x75, 0x18, 0x0F,
	0x22, 0x5F, 0x2A, 0x0F, 0x34, 0x5B, 0x5B, 0x28, 0x24, 0x20, 0x22, 0x11,
	0x28, 0x3F, 0x2C, 0x3D, 0x2A, 0x2C, 0x22, 0x15, 0x25, 0x1E, 0x2D, 0x14,
	0x10, 0x19, 0x3C, 0x12, 0x00, 0x04, 0x34, 0x09, 0x29, 0x26, 0x3B, 0x1C,
	0x07, 0x77, 0x5C, 0x02, 0x00, 0x01, 0x2E, 0x14, 0x55, 0x0F, 0x0F, 0x6D,
	0x26, 0x24, 0x1D, 0x11, 0x11, 0x28, 0x2A, 0x17, 0x3E, 0x36, 0x03, 0x22,
	0x0C, 0x5D, 0x00, 0x2E, 0x2F, 0x09, 0x5F, 0x73, 0x5A, 0x16, 0x5F, 0x2D,
	0x0C, 0x21, 0x14, 0x5F, 0x44, 0x1A, 0x01, 0x14, 0x34, 0x2F, 0x24, 0x1E,
	0x35, 0x05, 0x1B, 0x0E, 0x08, 0x56, 0x39, 0x28, 0x69, 0x06, 0x06, 0x23,
	0x5F, 0x12, 0x5B, 0x4E, 0x17, 0x12, 0x25, 0x02, 0x58, 0x2F, 0x40, 0x38,
	0x19, 0x29, 0x29, 0x5B, 0x29, 0x5C, 0x19, 0x08, 0x5E, 0x28, 0x07, 0x2A,
	0x2F, 0x58, 0x01, 0x07, 0x32, 0x1A, 0x5C, 0x32, 0x23, 0x53, 0x24, 0x3E,
	0x73, 0x5D, 0x12, 0x24, 0x0D, 0x71, 0x27, 0x26, 0x57, 0x18, 0x26, 0x24,
	0x0A, 0x5C, 0x21, 0x74, 0x1F, 0x0B, 0x56, 0x1F, 0x38, 0x39, 0x2E, 0x3C,
	0x3A, 0x15, 0x28, 0x4E, 0x59, 0x1D, 0x37, 0x5C, 0x13, 0x5F, 0x3B, 0x2E,
	0x05, 0x0B, 0x2D, 0x23, 0x15, 0x0A, 0x2E, 0x34, 0x1C, 0x72, 0x5A, 0x2C,
	0x3F, 0x11, 0x1B, 0x3B, 0x06, 0x17, 0x1F, 0x10, 0x28, 0x2A, 0x5A, 0x5D,
	0x38, 0x04, 0x29, 0x5B, 0x03, 0x2D, 0x3C, 0x19, 0x14, 0x5D, 0x26, 0x03,
	0x36, 0x1D, 0x0D, 0x0D, 0x36, 0x38, 0x1B, 0x33, 0x0A, 0x02, 0x06, 0x2D,
	0x09, 0x7A, 0x2A, 0x35, 0x00, 0x2A, 0x01, 0x2B, 0x0E, 0x5A, 0x20, 0x20,
	0x24, 0x34, 0x0F, 0x21, 0x2C, 0x3E, 0x3B, 0x29, 0x39, 0x04, 0x38, 0x25,
	0x05, 0x25, 0x74, 0x24, 0x22, 0x09, 0x23, 0x23, 0x5E, 0x0F, 0x08, 0x07,
	0x16, 0x36, 0x15, 0x2D, 0x3B, 0x0D, 0x0B, 0x03, 0x21, 0x00, 0x33, 0x5A,
	0x10, 0x14, 0x5B, 0x12, 0x23, 0x0E, 0x2B, 0x5B, 0x0D, 0x1E, 0x59, 0x20,
	0x3D, 0x1A, 0x25, 0x36, 0x2C, 0x5A, 0x3B, 0x2B, 0x02, 0x0D, 0x2F, 0x36,
	0x2E, 0x09, 0x04, 0x1C, 0x04, 0x54, 0x05, 0x41, 0x33, 0x74, 0x06, 0x0A,
	0x5A, 0x23, 0x2A, 0x15, 0x39, 0x25, 0x13, 0x0B, 0x14, 0x04, 0x1B, 0x3A,
	0x2C, 0x5F, 0x14, 0x2B, 0x29, 0x14, 0x2D, 0x20, 0x59, 0x0D, 0x15, 0x1A,
	0x54, 0x24, 0x52, 0x74, 0x3E, 0x29, 0x21, 0x0C, 0x2E, 0x1D, 0x1B, 0x29,
	0x3A, 0x28, 0x2A, 0x07, 0x02, 0x5E, 0x04, 0x5F, 0x55, 0x07, 0x59, 0x24,
	0x36, 0x15, 0x14, 0x53, 0x7B, 0x09, 0x58, 0x3E, 0x2A, 0x06, 0x1A, 0x17,
	0x25, 0x04, 0x0E, 0x0F, 0x34, 0x34, 0x1D, 0x21, 0x3E, 0x29, 0x0D, 0x0E,
	0x18, 0x5F, 0x00, 0x26, 0x04, 0x23, 0x1D, 0x31, 0x18, 0x5F, 0x73, 0x14,
	0x32, 0x2B, 0x58, 0x72, 0x54, 0x03, 0x57, 0x20, 0x6D, 0x19, 0x3B, 0x3B,
	0x5E, 0x2F, 0x47, 0x39, 0x0A, 0x26, 0x71, 0x1D, 0x0F, 0x34, 0x29, 0x06,
	0x2B, 0x50, 0x1E, 0x19, 0x24, 0x54, 0x00, 0x14, 0x32, 0x23, 0x00, 0x52,
	0x22, 0x0C, 0x09, 0x15, 0x52, 0x25, 0x40, 0x07, 0x47, 0x38, 0x1A, 0x0F,
	0x05, 0x3D, 0x28, 0x1F, 0x04, 0x16, 0x1C, 0x09, 0x22, 0x04, 0x03, 0x25,
	0x52, 0x3F, 0x33, 0x0A, 0x2F, 0x22, 0x37, 0x23, 0x75, 0x24, 0x32, 0x57,
	0x3F, 0x2B, 0x09, 0x07, 0x5C, 0x04, 0x71, 0x55, 0x4E, 0x27, 0x2F, 0x25,
	0x0E, 0x08, 0x20, 0x12, 0x0F, 0x3D, 0x57, 0x08, 0x2E, 0x2C, 0x21, 0x04,
	0x22, 0x25, 0x18, 0x19, 0x27, 0x20, 0x1C, 0x75, 0x01, 0x2C, 0x14, 0x23,
	0x0E, 0x08, 0x57, 0x1F, 0x2C, 0x04, 0x19, 0x57, 0x2A, 0x13, 0x28, 0x3F,
	0x19, 0x05, 0x3C, 0x16, 0x5C, 0x02, 0x2F, 0x09, 0x1B, 0x0F, 0x00, 0x18,
	0x08, 0x37, 0x20, 0x33, 0x3D, 0x03, 0x70, 0x09, 0x3B, 0x04, 0x3C, 0x0B,
	0x09, 0x30, 0x22, 0x0F, 0x33, 0x02, 0x2E, 0x2F, 0x22, 0x05, 0x18, 0x51,
	0x3A, 0x08, 0x18, 0x20, 0x11, 0x41, 0x3F, 0x0D, 0x1E, 0x0C, 0x27, 0x2C,
	0x12, 0x1B, 0x36, 0x18, 0x3F, 0x0F, 0x2F, 0x0B, 0x5C, 0x09, 0x34, 0x58,
	0x20, 0x03, 0x3D, 0x31, 0x06, 0x4E, 0x59, 0x04, 0x27, 0x14, 0x59, 0x07,
	0x1E, 0x2E, 0x03, 0x32, 0x24, 0x5D, 0x27, 0x20, 0x2D, 0x04, 0x33, 0x10,
	0x59, 0x13, 0x3B, 0x05, 0x35, 0x07, 0x17, 0x16, 0x18, 0x6D, 0x05, 0x23,
	0x18, 0x1F, 0x7A, 0x3E, 0x15, 0x04, 0x5D, 0x0A, 0x35, 0x2A, 0x5E, 0x04,
	0x16, 0x23, 0x30, 0x39, 0x0C, 0x27, 0x2B, 0x2B, 0x02, 0x1C, 0x6D, 0x0B,
	0x4E, 0x1B, 0x1F, 0x37, 0x24, 0x12, 0x14, 0x3C, 0x31, 0x5C, 0x3B, 0x5B,
	0x2F, 0x16, 0x58, 0x18, 0x36, 0x08, 0x24, 0x2E, 0x05, 0x20, 0x25, 0x36,
	0x2A, 0x22, 0x00, 0x3C, 0x06, 0x25, 0x36, 0x37, 0x2A, 0x20, 0x01, 0x12,
	0x2A, 0x04, 0x06, 0x5C, 0x4E, 0x16, 0x2F, 0x71, 0x20, 0x14, 0x2C, 0x25,
	0x14, 0x3A, 0x0F, 0x41, 0x08, 0x07, 0x5A, 0x03, 0x57, 0x2A, 0x0B, 0x18,
	0x2B, 0x5A, 0x3D, 0x15, 0x29, 0x34, 0x2B, 0x2F, 0x04, 0x2F, 0x34, 0x25,
	0x06, 0x28, 0x1E, 0x18, 0x2A, 0x07, 0x1A, 0x3D, 0x23, 0x28, 0x22, 0x76,
	0x1D, 0x00, 0x00, 0x2C, 0x05, 0x34, 0x30, 0x3F, 0x13, 0x23, 0x00, 0x35,
	0x3C, 0x39, 0x25, 0x3E, 0x2A, 0x1C, 0x38, 0x09, 0x06, 0x0C, 0x24, 0x27,
	0x15, 0x1F, 0x06, 0x16, 0x23, 0x0D, 0x1B, 0x06, 0x5A, 0x59, 0x70, 0x0F,
	0x12, 0x0F, 0x26, 0x76, 0x58, 0x55, 0x19, 0x5F, 0x73, 0x04, 0x0A, 0x26,
	0x3C, 0x72, 0x3E, 0x2F, 0x39, 0x06, 0x25, 0x20, 0x04, 0x2B, 0x06, 0x0E,
	0x25, 0x09, 0x0D, 0x1D, 0x2D, 0x3F, 0x08, 0x0B, 0x3A, 0x75, 0x07, 0x24,
	0x3B, 0x23, 0x32, 0x2E, 0x0C, 0x18, 0x52, 0x23, 0x0D, 0x54, 0x45, 0x00,
	0x74, 0x3D, 0x3B, 0x57, 0x5E, 0x6D, 0x1A, 0x4A, 0x14, 0x44, 0x0C, 0x55,
	0x31, 0x2F, 0x44, 0x0C, 0x47, 0x04, 0x5C, 0x11, 0x7B, 0x06, 0x56, 0x59,
	0x18, 0x34, 0x0E, 0x00, 0x0F, 0x40, 0x69, 0x55, 0x58, 0x1A, 0x19, 0x0A,
	0x02, 0x19, 0x08, 0x32, 0x72, 0x1F, 0x2B, 0x0D, 0x2D, 0x36, 0x05, 0x20,
	0x09, 0x3D, 0x12, 0x3D, 0x0C, 0x5F, 0x23, 0x0D, 0x25, 0x4E, 0x0D, 0x2F,
	0x33, 0x54, 0x19, 0x09, 0x52, 0x6D, 0x07, 0x24, 0x1A, 0x0F, 0x0A, 0x3E,
	0x4E, 0x18, 0x23, 0x0E, 0x1C, 0x35, 0x16, 0x06, 0x26, 0x1F, 0x09, 0x2C,
	0x3D, 0x72, 0x1F, 0x23, 0x36, 0x38, 0x3A, 0x09, 0x53, 0x21, 0x21, 0x0F,
	0x5B, 0x53, 0x0C, 0x01, 0x05, 0x04, 0x53, 0x3A, 0x2E, 0x2D, 0x26, 0x18,
	0x0F, 0x5A, 0x00, 0x22, 0x33, 0x1F, 0x24, 0x35, 0x54, 0x24, 0x00, 0x1B,
	0x0C, 0x09, 0x52, 0x45, 0x06, 0x0A, 0x16, 0x25, 0x23, 0x5B, 0x2E, 0x5C,
	0x54, 0x5F, 0x3B, 0x2F, 0x5E, 0x0F, 0x27, 0x53, 0x21, 0x27, 0x50, 0x03,
	0x13, 0x03, 0x1D, 0x58, 0x5A, 0x0C, 0x75, 0x03, 0x53, 0x57, 0x5E, 0x37,
	0x58, 0x02, 0x26, 0x29, 0x75, 0x21, 0x55, 0x57, 0x3E, 0x71, 0x59, 0x54,
	0x2B, 0x03, 0x73, 0x2E, 0x05, 0x58, 0x11, 0x00, 0x07, 0x30, 0x3B, 0x38,
	0x29, 0x2D, 0x2C, 0x21, 0x44, 0x1A, 0x21, 0x15, 0x3A, 0x0C, 0x0A, 0x55,
	0x52, 0x06, 0x06, 0x72, 0x24, 0x20, 0x01, 0x1E, 0x3B, 0x22, 0x12, 0x5C,
	0x11, 0x3B, 0x01, 0x56, 0x06, 0x3F, 0x75, 0x22, 0x27, 0x3E, 0x1D, 0x0D,
	0x06, 0x58, 0x07, 0x11, 0x09, 0x36, 0x0D, 0x00, 0x3A, 0x03, 0x36, 0x26,
	0x0D, 0x58, 0x77, 0x43, 0x17, 0x5A, 0x07, 0x0F, 0x27, 0x2A, 0x26, 0x06,
	0x30, 0x26, 0x2A, 0x3D, 0x08, 0x75, 0x3D, 0x05, 0x2F, 0x5D, 0x34, 0x19,
	0x3B, 0x5D, 0x0E, 0x16, 0x02, 0x2D, 0x45, 0x1B, 0x14, 0x05, 0x35, 0x0F,
	0x11, 0x69, 0x59, 0x2F, 0x23, 0x04, 0x03, 0x1B, 0x59, 0x5A, 0x44, 0x74,
	0x2A, 0x56, 0x14, 0x29, 0x72, 0x5B, 0x2E, 0x04, 0x44, 0x2C, 0x58, 0x4E,
	0x0C, 0x0E, 0x09, 0x54, 0x09, 0x17, 0x52, 0x70, 0x19, 0x11, 0x39, 0x21,
	0x77, 0x0A, 0x07, 0x3D, 0x06, 0x36, 0x58, 0x37, 0x5E, 0x20, 0x17, 0x2D,
	0x18, 0x16, 0x1A, 0x2D, 0x3B, 0x2D, 0x0D, 0x28, 0x01, 0x0D, 0x09, 0x26,
	0x0D, 0x36, 0x22, 0x02, 0x57, 0x1A, 0x76, 0x09, 0x51, 0x03, 0x5F, 0x3A,
	0x38, 0x03, 0x06, 0x33, 0x36, 0x15, 0x2E, 0x3D, 0x3F, 0x1A, 0x00, 0x20,
	0x1C, 0x2F, 0x75, 0x5A, 0x0F, 0x28, 0x5C, 0x32, 0x16, 0x16, 0x59, 0x28,
	0x0C, 0x0D, 0x59, 0x14, 0x38, 0x77, 0x01, 0x25, 0x20, 0x1D, 0x16, 0x2A,
	0x23, 0x41, 0x3F, 0x33, 0x34, 0x31, 0x0F, 0x5D, 0x20, 0x2A, 0x22, 0x22,
	0x0A, 0x26, 0x21, 0x28, 0x1A, 0x03, 0x35, 0x2B, 0x13, 0x5F, 0x5C, 0x00,
	0x3A, 0x58, 0x3E, 0x5D, 0x1A, 0x5B, 0x53, 0x56, 0x24, 0x01, 0x02, 0x53,
	0x58, 0x03, 0x2E, 0x54, 0x05, 0x39, 0x05, 0x6D, 0x1D, 0x18, 0x00, 0x52,
	0x31, 0x36, 0x56, 0x2D, 0x3D, 0x3A, 0x02, 0x58, 0x1C, 0x44, 0x74, 0x1B,
	0x2F, 0x2C, 0x5C, 0x30, 0x55, 0x4E, 0x04, 0x1A, 0x69, 0x20, 0x31, 0x16,
	0x3D, 0x75, 0x0A, 0x53, 0x24, 0x5A, 0x2B, 0x26, 0x13, 0x5D, 0x09, 0x73,
	0x1A, 0x56, 0x1F, 0x12, 0x12, 0x54, 0x29, 0x08, 0x5F, 0x23, 0x18, 0x52,
	0x45, 0x07, 0x7B, 0x55, 0x12, 0x28, 0x5E, 0x03, 0x3A, 0x56, 0x0F, 0x3B,
	0x35, 0x5A, 0x15, 0x02, 0x40, 0x09, 0x1C, 0x36, 0x08, 0x11, 0x15, 0x29,
	0x0D, 0x1C, 0x38, 0x1A, 0x35, 0x2F, 0x2D, 0x04, 0x08, 0x58, 0x08, 0x5F,
	0x0A, 0x34, 0x2B, 0x54, 0x3B, 0x05, 0x7A, 0x55, 0x27, 0x2C, 0x1B, 0x03,
	0x43, 0x04, 0x2B, 0x31, 0x03, 0x08, 0x09, 0x5D, 0x0E, 0x1B, 0x1C, 0x12,
	0x5C, 0x1D, 0x77, 0x34, 0x56, 0x22, 0x0E, 0x18, 0x0D, 0x54, 0x26, 0x00,
	0x38, 0x07, 0x32, 0x3D, 0x1F, 0x28, 0x06, 0x2B, 0x05, 0x5F, 0x3B, 0x29,
	0x12, 0x00, 0x0A, 0x36, 0x38, 0x0E, 0x22, 0x33, 0x00, 0x5A, 0x0E, 0x0C,
	0x02, 0x17, 0x3E, 0x02, 0x09, 0x11, 0x34, 0x23, 0x12, 0x1D, 0x06, 0x69,
	0x02, 0x12, 0x06, 0x28, 0x11, 0x26, 0x00, 0x1A, 0x00, 0x69, 0x39, 0x06,
	0x5C, 0x38, 0x33, 0x3B, 0x34, 0x1C, 0x19, 0x72, 0x20, 0x25, 0x3C, 0x2F,
	0x0B, 0x3F, 0x03, 0x03, 0x05, 0x6D, 0x38, 0x4A, 0x08, 0x0F, 0x00, 0x5C,
	0x14, 0x5B, 0x11, 0x69, 0x39, 0x32, 0x1B, 0x3C, 0x2D, 0x2D, 0x4E, 0x5D,
	0x1A, 0x2C, 0x18, 0x0E, 0x17, 0x09, 0x3A, 0x1F, 0x12, 0x20, 0x39, 0x2B,
	0x0F, 0x0A, 0x27, 0x5D, 0x71, 0x3B, 0x30, 0x2D, 0x25, 0x1A, 0x34, 0x14,
	0x0B, 0x0F, 0x28, 0x19, 0x2D, 0x57, 0x19, 0x37, 0x23, 0x28, 0x21, 0x0A,
	0x12, 0x27, 0x56, 0x58, 0x05, 0x3B, 0x5B, 0x27, 0x28, 0x11, 0x2C, 0x0A,
	0x17, 0x37, 0x27, 0x24, 0x09, 0x06, 0x22, 0x58, 0x76, 0x3A, 0x32, 0x5F,
	0x07, 0x05, 0x3E, 0x10, 0x59, 0x3C, 0x72, 0x01, 0x0D, 0x2F, 0x01, 0x0D,
	0x22, 0x31, 0x3C, 0x3F, 0x24, 0x04, 0x34, 0x0F, 0x27, 0x18, 0x1C, 0x32,
	0x02, 0x02, 0x20, 0x1C, 0x56, 0x2D, 0x31, 0x15, 0x5F, 0x35, 0x09, 0x32,
	0x38, 0x3A, 0x55, 0x1D, 0x1F, 0x09, 0x15, 0x10, 0x18, 0x1D, 0x0B, 0x21,
	0x33, 0x04, 0x0D, 0x73, 0x0A, 0x36, 0x01, 0x2E, 0x7B, 0x34, 0x32, 0x5B,
	0x5D, 0x21, 0x1F, 0x0D, 0x0B, 0x2E, 0x08, 0x19, 0x38, 0x39, 0x29, 0x27,
	0x06, 0x36, 0x09, 0x5A, 0x29, 0x3C, 0x0D, 0x56, 0x0D, 0x29, 0x1A, 0x54,
	0x0A, 0x5B, 0x77, 0x43, 0x1B, 0x1A, 0x09, 0x75, 0x55, 0x39, 0x5D, 0x06,
	0x16, 0x38, 0x22, 0x14, 0x53, 0x29, 0x59, 0x15, 0x0B, 0x5F, 0x03, 0x3B,
	0x18, 0x26, 0x5F, 0x0E, 0x1A, 0x25, 0x21, 0x1D, 0x3B, 0x43, 0x35, 0x02,
	0x08, 0x01, 0x05, 0x22, 0x25, 0x2D, 0x23, 0x28, 0x03, 0x03, 0x52, 0x13,
	0x28, 0x18, 0x17, 0x07, 0x16, 0x20, 0x1B, 0x56, 0x2A, 0x0C, 0x00, 0x02,
	0x0A, 0x0A, 0x1A, 0x3E, 0x34, 0x18, 0x03, 0x0E, 0x28, 0x4A, 0x06, 0x2C,
	0x1A, 0x1C, 0x4A, 0x02, 0x22, 0x75, 0x0F, 0x15, 0x18, 0x3D, 0x69, 0x43,
	0x04, 0x2D, 0x1F, 0x16, 0x09, 0x38, 0x2D, 0x1F, 0x21, 0x38, 0x3B, 0x2F,
	0x18, 0x2F, 0x1D, 0x13, 0x04, 0x3F, 0x0E, 0x5B, 0x04, 0x19, 0x03, 0x16,
	0x22, 0x58, 0x18, 0x22, 0x15, 0x20, 0x2D, 0x58, 0x2A, 0x26, 0x1C, 0x3B,
	0x39, 0x3E, 0x13, 0x43, 0x2D, 0x39, 0x3A, 0x70, 0x47, 0x02, 0x19, 0x0C,
	0x24, 0x3F, 0x37, 0x17, 0x11, 0x23, 0x2E, 0x4A, 0x45, 0x13, 0x71, 0x5D,
	0x59, 0x58, 0x08, 0x16, 0x55, 0x58, 0x06, 0x5C, 0x73, 0x2D, 0x59, 0x2F,
	0x5B, 0x73, 0x5C, 0x32, 0x58, 0x1F, 0x32, 0x0D, 0x00, 0x18, 0x1B, 0x75,
	0x1F, 0x35, 0x38, 0x3C, 0x12, 0x05, 0x51, 0x37, 0x32, 0x34, 0x0A, 0x57,
	0x01, 0x23, 0x34, 0x39, 0x08, 0x1D, 0x00, 0x35, 0x47, 0x20, 0x09, 0x1B,
	0x31, 0x09, 0x31, 0x06, 0x11, 0x0E, 0x02, 0x58, 0x0C, 0x3E, 0x2A, 0x59,
	0x04, 0x2C, 0x33, 0x04, 0x3B, 0x0E, 0x26, 0x3B, 0x2C, 0x02, 0x08, 0x1D,
	0x18, 0x2B, 0x07, 0x34, 0x5A, 0x5A, 0x74, 0x27, 0x02, 0x0F, 0x04, 0x2D,
	0x43, 0x18, 0x2A, 0x04, 0x10, 0x14, 0x32, 0x00, 0x23, 0x0D, 0x02, 0x10,
	0x38, 0x5A, 0x0A, 0x3E, 0x31, 0x0B, 0x0F, 0x06, 0x3C, 0x3B, 0x3C, 0x01,
	0x03, 0x5C, 0x57, 0x26, 0x1B, 0x3B, 0x3D, 0x32, 0x57, 0x21, 0x0C, 0x01,
	0x0F, 0x37, 0x40, 0x28, 0x05, 0x00, 0x37, 0x5D, 0x2C, 0x5E, 0x27, 0x1C,
	0x12, 0x33, 0x43, 0x09, 0x29, 0x0D, 0x3B, 0x3F, 0x35, 0x25, 0x3E, 0x17,
	0x36, 0x28, 0x19, 0x1C, 0x20, 0x01, 0x2E, 0x1E, 0x33, 0x28, 0x43, 0x0D,
	0x03, 0x20, 0x2F, 0x1C, 0x59, 0x59, 0x0A, 0x25, 0x14, 0x04, 0x17, 0x3A,
	0x18, 0x18, 0x2F, 0x0D, 0x0E, 0x00, 0x2F, 0x00, 0x3A, 0x31, 0x27, 0x2D,
	0x23, 0x07, 0x21, 0x03, 0x09, 0x15, 0x0A, 0x3C, 0x31, 0x24, 0x11, 0x2A,
	0x20, 0x76, 0x01, 0x2A, 0x03, 0x27, 0x2F, 0x0F, 0x36, 0x16, 0x07, 0x73,
	0x27, 0x38, 0x3D, 0x5C, 0x15, 0x04, 0x13, 0x16, 0x19, 0x34, 0x2D, 0x08,
	0x0F, 0x12, 0x34, 0x5A, 0x54, 0x2B, 0x31, 0x12, 0x2A, 0x51, 0x05, 0x02,
	0x69, 0x18, 0x3B, 0x19, 0x12, 0x26, 0x00, 0x2F, 0x2B, 0x07, 0x74, 0x19,
	0x0F, 0x3C, 0x52, 0x1B, 0x0F, 0x09, 0x05, 0x5D, 0x76, 0x2D, 0x22, 0x5B,
	0x09, 0x2F, 0x5E, 0x25, 0x01, 0x3C, 0x0E, 0x26, 0x54, 0x57, 0x27, 0x75,
	0x39, 0x39, 0x5F, 0x58, 0x3B, 0x3F, 0x37, 0x3E, 0x02, 0x10, 0x29, 0x15,
	0x5D, 0x3E, 0x24, 0x15, 0x10, 0x56, 0x3D, 0x72, 0x35, 0x55, 0x00, 0x0E,
	0x11, 0x28, 0x0F, 0x0A, 0x5E, 0x75, 0x29, 0x2D, 0x5D, 0x1F, 0x06, 0x5A,
	0x14, 0x1D, 0x3D, 0x72, 0x54, 0x25, 0x14, 0x3C, 0x07, 0x08, 0x52, 0x45,
	0x38, 0x16, 0x43, 0x4E, 0x28, 0x3F, 0x10, 0x54, 0x1B, 0x18, 0x58, 0x38,
	0x0D, 0x37, 0x26, 0x3A, 0x20, 0x5A, 0x10, 0x57, 0x01, 0x72, 0x59, 0x0A,
	0x2A, 0x3B, 0x05, 0x0E, 0x0D, 0x1A, 0x44, 0x0A, 0x2A, 0x10, 0x39, 0x33,
	0x05, 0x38, 0x29, 0x29, 0x5C, 0x2F, 0x1B, 0x36, 0x19, 0x12, 0x2F, 0x1E,
	0x30, 0x3A, 0x33, 0x0C, 0x01, 0x00, 0x0D, 0x5D, 0x3A, 0x35, 0x50, 0x06,
	0x1D, 0x72, 0x07, 0x04, 0x16, 0x1E, 0x18, 0x0F, 0x0F, 0x58, 0x3F, 0x33,
	0x28, 0x0E, 0x23, 0x0A, 0x03, 0x1A, 0x23, 0x26, 0x09, 0x21, 0x38, 0x05,
	0x22, 0x09, 0x70, 0x22, 0x22, 0x1A, 0x2E, 0x24, 0x0F, 0x59, 0x05, 0x3C,
	0x76, 0x3C, 0x2C, 0x24, 0x0F, 0x07, 0x55, 0x50, 0x2C, 0x02, 0x25, 0x2D,
	0x34, 0x21, 0x25, 0x16, 0x54, 0x25, 0x1C, 0x19, 0x16, 0x0F, 0x2F, 0x3F,
	0x12, 0x15, 0x1B, 0x33, 0x1F, 0x52, 0x77, 0x20, 0x19, 0x0B, 0x59, 0x0E,
	0x1B, 0x04, 0x17, 0x3F, 0x73, 0x38, 0x04, 0x3C, 0x00, 0x7A, 0x3E, 0x56,
	0x1D, 0x1D, 0x15, 0x3E, 0x53, 0x3A, 0x44, 0x37, 0x1A, 0x39, 0x1A, 0x21,
	0x0A, 0x1E, 0x13, 0x05, 0x07, 0x2F, 0x06, 0x2E, 0x1E, 0x05, 0x36, 0x3E,
	0x56, 0x24, 0x27, 0x77, 0x24, 0x30, 0x3D, 0x5A, 0x0D, 0x24, 0x2F, 0x1A,
	0x5A, 0x06, 0x16, 0x2A, 0x3A, 0x0E, 0x1B, 0x05, 0x14, 0x3C, 0x1D, 0x25,
	0x09, 0x29, 0x5C, 0x21, 0x0D, 0x34, 0x00, 0x2D, 0x3F, 0x2F, 0x27, 0x53,
	0x24, 0x1F, 0x07, 0x0F, 0x55, 0x38, 0x5D, 0x15, 0x5D, 0x1B, 0x39, 0x5F,
	0x71, 0x22, 0x02, 0x17, 0x2E, 0x3B, 0x43, 0x10, 0x2C, 0x22, 0x1A, 0x00,
	0x0E, 0x0B, 0x2C, 0x11, 0x0A, 0x18, 0x37, 0x5C, 0x76, 0x14, 0x52, 0x2B,
	0x18, 0x69, 0x20, 0x18, 0x5A, 0x01, 0x11, 0x43, 0x00, 0x3B, 0x5B, 0x0D,
	0x5E, 0x4A, 0x3B, 0x44, 0x13, 0x0D, 0x07, 0x26, 0x1B, 0x74, 0x5B, 0x57,
	0x1C, 0x0E, 0x74, 0x38, 0x58, 0x3C, 0x1A, 0x00, 0x43, 0x27, 0x41, 0x52,
	0x28, 0x1A, 0x22, 0x1E, 0x18, 0x33, 0x19, 0x02, 0x41, 0x04, 0x2F, 0x1E,
	0x27, 0x1E, 0x3B, 0x04, 0x26, 0x3B, 0x58, 0x00, 0x05, 0x0A, 0x07, 0x5A,
	0x22, 0x2C, 0x5E, 0x52, 0x0C, 0x3E, 0x2E, 0x1D, 0x03, 0x20, 0x3C, 0x69,
	0x47, 0x16, 0x18, 0x0A, 0x10, 0x0E, 0x15, 0x1C, 0x18, 0x20, 0x5A, 0x2D,
	0x5B, 0x1B, 0x7A, 0x5A, 0x09, 0x58, 0x32, 0x29, 0x34, 0x53, 0x20, 0x12,
	0x74, 0x28, 0x54, 0x22, 0x3F, 0x14, 0x00, 0x2B, 0x03, 0x59, 0x25, 0x34,
	0x4E, 0x5F, 0x09, 0x24, 0x3E, 0x2B, 0x18, 0x27, 0x7B, 0x00, 0x53, 0x21,
	0x27, 0x11, 0x27, 0x31, 0x0D, 0x04, 0x04, 0x2A, 0x14, 0x21, 0x52, 0x3B,
	0x5C, 0x04, 0x27, 0x29, 0x69, 0x15, 0x55, 0x26, 0x2D, 0x28, 0x2A, 0x2D,
	0x07, 0x19, 0x31, 0x2B, 0x56, 0x22, 0x1E, 0x0F, 0x43, 0x16, 0x00, 0x5C,
	0x2B, 0x09, 0x31, 0x5D, 0x44, 0x75, 0x47, 0x18, 0x00, 0x58, 0x25, 0x2A,
	0x0B, 0x5C, 0x3B, 0x21, 0x05, 0x4E, 0x1D, 0x1F, 0x74, 0x14, 0x07, 0x28,
	0x1F, 0x2E, 0x0E, 0x36, 0x22, 0x04, 0x30, 0x1A, 0x15, 0x14, 0x1C, 0x17,
	0x28, 0x58, 0x3C, 0x06, 0x74, 0x0A, 0x12, 0x1A, 0x58, 0x15, 0x5D, 0x12,
	0x41, 0x40, 0x35, 0x19, 0x10, 0x1F, 0x05, 0x0F, 0x01, 0x19, 0x08, 0x04,
	0x2A, 0x5F, 0x15, 0x00, 0x5F, 0x38, 0x00, 0x58, 0x5E, 0x11, 0x17, 0x20,
	0x36, 0x2F, 0x24, 0x24, 0x35, 0x2E, 0x1C, 0x09, 0x15, 0x3A, 0x00, 0x1D,
	0x21, 0x0D, 0x14, 0x2F, 0x26, 0x5B, 0x0B, 0x43, 0x15, 0x28, 0x3C, 0x2A,
	0x58, 0x1B, 0x0A, 0x08, 0x08, 0x34, 0x06, 0x36, 0x01, 0x21, 0x0F, 0x05,
	0x03, 0x1C, 0x70, 0x3D, 0x17, 0x05, 0x31, 0x2C, 0x0E, 0x0C, 0x2D, 0x2E,
	0x13, 0x25, 0x13, 0x02, 0x0A, 0x7B, 0x02, 0x0E, 0x38, 0x5E, 0x70, 0x24,
	0x03, 0x03, 0x3F, 0x0E, 0x15, 0x30, 0x02, 0x1F, 0x38, 0x1A, 0x27, 0x2F,
	0x00, 0x2D, 0x2A, 0x14, 0x39, 0x21, 0x12, 0x1D, 0x23, 0x08, 0x5B, 0x24,
	0x59, 0x2D, 0x3E, 0x07, 0x72, 0x08, 0x0B, 0x2F, 0x40, 0x10, 0x07, 0x04,
	0x1B, 0x0A, 0x75, 0x1F, 0x16, 0x37, 0x5F, 0x0A, 0x47, 0x09, 0x34, 0x0A,
	0x18, 0x21, 0x0F, 0x0C, 0x1F, 0x23, 0x3A, 0x51, 0x05, 0x06, 0x24, 0x1D,
	0x2B, 0x19, 0x1F, 0x08, 0x06, 0x59, 0x5C, 0x23, 0x2E, 0x2A, 0x33, 0x06,
	0x2A, 0x2D, 0x01, 0x19, 0x0A, 0x0C, 0x2A, 0x3F, 0x17, 0x59, 0x40, 0x21,
	0x14, 0x27, 0x04, 0x11, 0x13, 0x04, 0x2B, 0x04, 0x09, 0x3B, 0x16, 0x12,
	0x28, 0x59, 0x0F, 0x04, 0x0A, 0x17, 0x5C, 0x05, 0x3B, 0x0A, 0x17, 0x18,
	0x13, 0x55, 0x31, 0x25, 0x0E, 0x7A, 0x5B, 0x00, 0x09, 0x3C, 0x0E, 0x21,
	0x23, 0x28, 0x0C, 0x75, 0x1B, 0x23, 0x34, 0x0A, 0x0A, 0x16, 0x00, 0x08,
	0x18, 0x69, 0x28, 0x00, 0x1D, 0x19, 0x34, 0x1C, 0x58, 0x3F, 0x06, 0x1B,
	0x29, 0x00, 0x01, 0x06, 0x0C, 0x2E, 0x29, 0x22, 0x06, 0x1A, 0x58, 0x52,
	0x36, 0x1B, 0x06, 0x2D, 0x38, 0x1B, 0x5A, 0x2D, 0x2A, 0x05, 0x04, 0x06,
	0x2D, 0x2B, 0x10, 0x28, 0x06, 0x14, 0x1C, 0x51, 0x28, 0x5B, 0x3A, 0x0E,
	0x15, 0x3D, 0x5B, 0x35, 0x06, 0x37, 0x0A, 0x23, 0x6D, 0x2D, 0x15, 0x1F,
	0x2C, 0x69, 0x36, 0x0A, 0x22, 0x40, 0x05, 0x3B, 0x51, 0x17, 0x5E, 0x6D,
	0x36, 0x15, 0x57, 0x52, 0x37, 0x26, 0x04, 0x28, 0x3C, 0x23, 0x18, 0x23,
	0x45, 0x5A, 0x32, 0x1E, 0x23, 0x57, 0x18, 0x71, 0x47, 0x25, 0x08, 0x2E,
	0x14, 0x58, 0x4A, 0x1B, 0x3A, 0x0A, 0x09, 0x19, 0x1D, 0x3F, 0x70, 0x06,
	0x0F, 0x08, 0x0E, 0x10, 0x55, 0x29, 0x56, 0x26, 0x38, 0x3B, 0x57, 0x38,
	0x38, 0x17, 0x1A, 0x4A, 0x2C, 0x28, 0x33, 0x14, 0x07, 0x5E, 0x0A, 0x23,
	0x1C, 0x2F, 0x3D, 0x00, 0x17, 0x0F, 0x08, 0x17, 0x25, 0x0B, 0x01, 0x3B,
	0x0C, 0x3D, 0x0A, 0x14, 0x0F, 0x23, 0x00, 0x06, 0x55, 0x0E, 0x1A, 0x12,
	0x29, 0x54, 0x4A, 0x5F, 0x33, 0x38, 0x38, 0x06, 0x17, 0x0C, 0x37, 0x54,
	0x52, 0x45, 0x40, 0x15, 0x04, 0x35, 0x57, 0x5A, 0x34, 0x55, 0x4E, 0x41,
	0x18, 0x28, 0x54, 0x32, 0x17, 0x08, 0x12, 0x55, 0x24, 0x08, 0x3C, 0x70,
	0x47, 0x57, 0x02, 0x1B, 0x0E, 0x1E, 0x08, 0x3E, 0x06, 0x2D, 0x35, 0x50,
	0x0D, 0x1E, 0x1B, 0x1F, 0x2C, 0x09, 0x3E, 0x6D, 0x0B, 0x33, 0x38, 0x3E,
	0x21, 0x06, 0x13, 0x16, 0x3B, 0x03, 0x09, 0x0A, 0x1E, 0x52, 0x3A, 0x3F,
	0x55, 0x58, 0x0C, 0x24, 0x04, 0x27, 0x36, 0x5A, 0x18, 0x14, 0x4A, 0x1F,
	0x40, 0x14, 0x1A, 0x30, 0x34, 0x2D, 0x20, 0x0F, 0x0C, 0x28, 0x0A, 0x73,
	0x1E, 0x04, 0x14, 0x59, 0x2B, 0x01, 0x34, 0x2D, 0x21, 0x12, 0x26, 0x11,
	0x3A, 0x11, 0x16, 0x1D, 0x50, 0x39, 0x31, 0x15, 0x55, 0x27, 0x19, 0x02,
	0x30, 0x18, 0x10, 0x29, 0x3D, 0x2C, 0x39, 0x0A, 0x1A, 0x44, 0x00, 0x43,
	0x52, 0x2D, 0x2D, 0x18, 0x08, 0x34, 0x07, 0x18, 0x6D, 0x05, 0x17, 0x03,
	0x0A, 0x18, 0x21, 0x05, 0x3F, 0x1D, 0x03, 0x43, 0x23, 0x3A, 0x5A, 0x00,
	0x3D, 0x02, 0x07, 0x24, 0x69, 0x22, 0x59, 0x38, 0x44, 0x0A, 0x03, 0x30,
	0x2C, 0x07, 0x26, 0x3A, 0x58, 0x0F, 0x2A, 0x75, 0x1D, 0x36, 0x57, 0x08,
	0x35, 0x3F, 0x2C, 0x34, 0x19, 0x31, 0x03, 0x07, 0x23, 0x28, 0x2E, 0x14,
	0x37, 0x3A, 0x3D, 0x37, 0x03, 0x35, 0x14, 0x3A, 0x2D, 0x47, 0x4E, 0x3E,
	0x2F, 0x0F, 0x04, 0x39, 0x07, 0x04, 0x7A, 0x08, 0x06, 0x5A, 0x01, 0x2E,
	0x2F, 0x18, 0x3F, 0x18, 0x72, 0x20, 0x26, 0x56, 0x58, 0x18, 0x09, 0x30,
	0x1A, 0x5A, 0x6D, 0x43, 0x04, 0x20, 0x5D, 0x74, 0x07, 0x16, 0x0C, 0x00,
	0x20, 0x34, 0x32, 0x04, 0x3C, 0x12, 0x5C, 0x54, 0x2C, 0x01, 0x1A, 0x5C,
	0x54, 0x45, 0x5B, 0x25, 0x59, 0x2A, 0x5E, 0x3D, 0x37, 0x1A, 0x30, 0x24,
	0x09, 0x13, 0x3E, 0x3B, 0x1A, 0x5E, 0x37, 0x05, 0x3B, 0x06, 0x3B, 0x28,
	0x5D, 0x38, 0x5E, 0x5B, 0x01, 0x5B, 0x52, 0x08, 0x21, 0x6D, 0x00, 0x17,
	0x56, 0x3E, 0x2E, 0x08, 0x14, 0x41, 0x3C, 0x28, 0x2A, 0x57, 0x20, 0x2F,
	0x2F, 0x29, 0x36, 0x1D, 0x27, 0x38, 0x07, 0x38, 0x14, 0x0D, 0x2F, 0x15,
	0x09, 0x29, 0x5F, 0x26, 0x35, 0x00, 0x0D, 0x03, 0x0A, 0x01, 0x0E, 0x2D,
	0x5C, 0x2B, 0x00, 0x27, 0x59, 0x3F, 0x34, 0x02, 0x0F, 0x5D, 0x0E, 0x18,
	0x28, 0x31, 0x58, 0x28, 0x36, 0x15, 0x10, 0x45, 0x44, 0x29, 0x24, 0x19,
	0x41, 0x24, 0x06, 0x18, 0x2E, 0x28, 0x59, 0x15, 0x59, 0x0D, 0x36, 0x1F,
	0x71, 0x1A, 0x25, 0x59, 0x5E, 0x18, 0x01, 0x37, 0x04, 0x52, 0x1A, 0x04,
	0x0D, 0x56, 0x1E, 0x0C, 0x5B, 0x14, 0x3C, 0x5C, 0x1A, 0x02, 0x39, 0x22,
	0x5F, 0x7A, 0x25, 0x04, 0x0F, 0x29, 0x73, 0x24, 0x27, 0x59, 0x3D, 0x1A,
	0x2A, 0x13, 0x22, 0x0D, 0x3A, 0x5E, 0x15, 0x07, 0x26, 0x76, 0x38, 0x17,
	0x3B, 0x31, 0x77, 0x58, 0x27, 0x1C, 0x2A, 0x37, 0x1D, 0x05, 0x5D, 0x5F,
	0x12, 0x08, 0x0F, 0x5F, 0x44, 0x76, 0x36, 0x51, 0x5A, 0x02, 0x26, 0x5E,
	0x51, 0x20, 0x09, 0x2D, 0x55, 0x20, 0x1F, 0x20, 0x7B, 0x16, 0x28, 0x09,
	0x1F, 0x13, 0x1F, 0x15, 0x03, 0x33, 0x0F, 0x01, 0x16, 0x37, 0x0E, 0x73,
	0x01, 0x00, 0x19, 0x58, 0x16, 0x22, 0x18, 0x2C, 0x12, 0x34, 0x28, 0x2C,
	0x27, 0x3C, 0x3A, 0x5C, 0x34, 0x26, 0x08, 0x10, 0x3D, 0x35, 0x37, 0x38,
	0x36, 0x26, 0x2E, 0x3C, 0x31, 0x05, 0x35, 0x37, 0x16, 0x05, 0x37, 0x0A,
	0x06, 0x1D, 0x53, 0x17, 0x3D, 0x4E, 0x2C, 0x5F, 0x15, 0x07, 0x0B, 0x1C,
	0x40, 0x11, 0x55, 0x2E, 0x19, 0x3F, 0x26, 0x1C, 0x53, 0x26, 0x29, 0x33,
	0x5C, 0x53, 0x36, 0x3A, 0x1B, 0x58, 0x52, 0x1D, 0x0A, 0x7B, 0x54, 0x4A,
	0x06, 0x40, 0x2E, 0x39, 0x38, 0x41, 0x5E, 0x03, 0x1A, 0x59, 0x14, 0x3E,
	0x09, 0x16, 0x26, 0x36, 0x13, 0x08, 0x18, 0x11, 0x14, 0x33, 0x3A, 0x55,
	0x53, 0x41, 0x44, 0x35, 0x27, 0x32, 0x24, 0x0E, 0x31, 0x0B, 0x53, 0x45,
	0x33, 0x12, 0x5C, 0x55, 0x1A, 0x3B, 0x70, 0x47, 0x34, 0x5C, 0x13, 0x0A,
	0x5C, 0x54, 0x5D, 0x44, 0x0E, 0x1E, 0x2F, 0x5E, 0x0D, 0x12, 0x47, 0x29,
	0x1B, 0x21, 0x69, 0x20, 0x14, 0x5B, 0x53, 0x1A, 0x0D, 0x2D, 0x5C, 0x03,
	0x15, 0x07, 0x03, 0x1C, 0x11, 0x74, 0x02, 0x32, 0x08, 0x25, 0x30, 0x1F,
	0x32, 0x56, 0x25, 0x04, 0x16, 0x27, 0x5C, 0x18, 0x35, 0x43, 0x00, 0x45,
	0x2C, 0x7B, 0x1A, 0x0E, 0x03, 0x5F, 0x3B, 0x26, 0x29, 0x3D, 0x2D, 0x05,
	0x21, 0x13, 0x2A, 0x52, 0x01, 0x20, 0x58, 0x24, 0x1E, 0x32, 0x5C, 0x0A,
	0x5E, 0x3E, 0x13, 0x3E, 0x18, 0x00, 0x32, 0x14, 0x21, 0x16, 0x0D, 0x20,
	0x38, 0x05, 0x07, 0x0C, 0x03, 0x09, 0x38, 0x54, 0x21, 0x2D, 0x32, 0x29,
	0x54, 0x09, 0x53, 0x1B, 0x20, 0x07, 0x5A, 0x3F, 0x3B, 0x47, 0x35, 0x14,
	0x25, 0x00, 0x1E, 0x0C, 0x08, 0x23, 0x7A, 0x1A, 0x56, 0x3C, 0x3D, 0x69,
	0x09, 0x36, 0x57, 0x53, 0x30, 0x43, 0x23, 0x5C, 0x29, 0x21, 0x1C, 0x56,
	0x24, 0x12, 0x34, 0x1A, 0x36, 0x03, 0x12, 0x31, 0x14, 0x14, 0x38, 0x5F,
	0x2A, 0x26, 0x56, 0x25, 0x07, 0x12, 0x21, 0x06, 0x08, 0x22, 0x71, 0x2B,
	0x56, 0x58, 0x00, 0x18, 0x2B, 0x35, 0x09, 0x31, 0x1A, 0x16, 0x15, 0x37,
	0x3D, 0x69, 0x26, 0x11, 0x24, 0x22, 0x26, 0x04, 0x39, 0x23, 0x5F, 0x7A,
	0x23, 0x33, 0x06, 0x0D, 0x6D, 0x2F, 0x05, 0x2A, 0x52, 0x75, 0x05, 0x06,
	0x3A, 0x24, 0x70, 0x2D, 0x20, 0x23, 0x58, 0x18, 0x38, 0x32, 0x0B, 0x5E,
	0x73, 0x5C, 0x28, 0x19, 0x2F, 0x30, 0x3A, 0x00, 0x58, 0x44, 0x24, 0x5C,
	0x06, 0x38, 0x5B, 0x36, 0x54, 0x28, 0x29, 0x5C, 0x7A, 0x2D, 0x31, 0x38,
	0x58, 0x38, 0x22, 0x09, 0x1A, 0x1B, 0x14, 0x59, 0x12, 0x08, 0x09, 0x2C,
	0x00, 0x2D, 0x2D, 0x08, 0x37, 0x0A, 0x15, 0x14, 0x2D, 0x2E, 0x1B, 0x2F,
	0x21, 0x31, 0x0D, 0x05, 0x00, 0x20, 0x5A, 0x77, 0x21, 0x27, 0x1B, 0x5C,
	0x74, 0x3E, 0x30, 0x57, 0x33, 0x09, 0x38, 0x2F, 0x01, 0x22, 0x27, 0x1A,
	0x12, 0x59, 0x3C, 0x33, 0x24, 0x4A, 0x04, 0x03, 0x0B, 0x19, 0x50, 0x5D,
	0x09, 0x05, 0x3F, 0x55, 0x2D, 0x58, 0x2C, 0x3A, 0x22, 0x27, 0x05, 0x75,
	0x1C, 0x19, 0x58, 0x52, 0x0C, 0x58, 0x0F, 0x21, 0x32, 0x08, 0x3F, 0x09,
	0x3F, 0x3C, 0x29, 0x5D, 0x14, 0x57, 0x31, 0x74, 0x23, 0x19, 0x37, 0x1E,
	0x77, 0x5D, 0x27, 0x17, 0x38, 0x24, 0x34, 0x0F, 0x5D, 0x53, 0x1B, 0x19,
	0x20, 0x18, 0x19, 0x03, 0x20, 0x59, 0x3C, 0x06, 0x26, 0x36, 0x52, 0x59,
	0x5F, 0x27, 0x2A, 0x1B, 0x17, 0x2C, 0x0A, 0x02, 0x56, 0x1C, 0x3B, 0x37,
	0x20, 0x50, 0x19, 0x06, 0x15, 0x1F, 0x15, 0x17, 0x3B, 0x23, 0x20, 0x50,
	0x5E, 0x0F, 0x3A, 0x05, 0x32, 0x08, 0x5E, 0x1B, 0x43, 0x0D, 0x3D, 0x1A,
	0x75, 0x29, 0x29, 0x3C, 0x52, 0x7B, 0x2D, 0x0B, 0x59, 0x1B, 0x0B, 0x16,
	0x28, 0x2B, 0x24, 0x34, 0x1B, 0x27, 0x03, 0x28, 0x0F, 0x19, 0x0D, 0x18,
	0x53, 0x7B, 0x2F, 0x02, 0x1A, 0x1F, 0x37, 0x18, 0x31, 0x26, 0x25, 0x09,
	0x03, 0x2A, 0x18, 0x0D, 0x16, 0x35, 0x39, 0x45, 0x24, 0x71, 0x0D, 0x0D,
	0x28, 0x3A, 0x2F, 0x3E, 0x28, 0x00, 0x40, 0x23, 0x3B, 0x54, 0x03, 0x2A,
	0x36, 0x16, 0x2C, 0x34, 0x09, 0x2E, 0x26, 0x18, 0x1C, 0x0E, 0x11, 0x14,
	0x23, 0x2B, 0x33, 0x73, 0x3E, 0x10, 0x1E, 0x26, 0x13, 0x3D, 0x0E, 0x0B,
	0x26, 0x0D, 0x20, 0x0D, 0x2F, 0x3F, 0x05, 0x1A, 0x28, 0x56, 0x20, 0x2D,
	0x2A, 0x18, 0x2F, 0x1B, 0x21, 0x38, 0x19, 0x45, 0x08, 0x38, 0x14, 0x58,
	0x1D, 0x5A, 0x1A, 0x15, 0x03, 0x02, 0x00, 0x70, 0x35, 0x27, 0x5F, 0x23,
	0x09, 0x06, 0x26, 0x24, 0x3A, 0x0E, 0x3F, 0x2B, 0x1C, 0x22, 0x2F, 0x1F,
	0x0B, 0x39, 0x01, 0x16, 0x5B, 0x27, 0x5D, 0x2E, 0x6D, 0x23, 0x15, 0x27,
	0x27, 0x17, 0x5D, 0x38, 0x58, 0x5E, 0x0E, 0x3D, 0x08, 0x03, 0x0F, 0x74,
	0x54, 0x15, 0x18, 0x00, 0x13, 0x16, 0x27, 0x0C, 0x04, 0x6D, 0x25, 0x19,
	0x3F, 0x05, 0x35, 0x05, 0x59, 0x38, 0x08, 0x17, 0x2B, 0x18, 0x38, 0x09,
	0x2D, 0x36, 0x0A, 0x36, 0x5F, 0x3B, 0x1B, 0x22, 0x0D, 0x1E, 0x36, 0x5F,
	0x2B, 0x01, 0x5B, 0x07, 0x2E, 0x39, 0x2D, 0x5F, 0x2F, 0x5D, 0x53, 0x1D,
	0x05, 0x0C, 0x09, 0x14, 0x0B, 0x5F, 0x18, 0x3F, 0x13, 0x41, 0x24, 0x38,
	0x0D, 0x2C, 0x24, 0x3E, 0x0B, 0x5F, 0x19, 0x3D, 0x20, 0x74, 0x24, 0x23,
	0x37, 0x31, 0x7B, 0x35, 0x09, 0x36, 0x5D, 0x1A, 0x34, 0x05, 0x5B, 0x07,
	0x23, 0x3D, 0x00, 0x5C, 0x44, 0x17, 0x36, 0x29, 0x28, 0x02, 0x10, 0x59,
	0x2F, 0x58, 0x03, 0x24, 0x3A, 0x50, 0x23, 0x5E, 0x25, 0x01, 0x27, 0x04,
	0x1D, 0x73, 0x0D, 0x26, 0x02, 0x58, 0x16, 0x20, 0x52, 0x08, 0x0C, 0x26,
	0x1A, 0x28, 0x41, 0x2E, 0x75, 0x04, 0x38, 0x07, 0x53, 0x25, 0x35, 0x57,
	0x5F, 0x32, 0x24, 0x23, 0x3B, 0x1D, 0x00, 0x10, 0x20, 0x23, 0x5A, 0x05,
	0x00, 0x15, 0x39, 0x58, 0x32, 0x35, 0x22, 0x50, 0x1D, 0x20, 0x3B, 0x5B,
	0x05, 0x20, 0x5E, 0x0C, 0x3F, 0x51, 0x22, 0x27, 0x38, 0x25, 0x31, 0x3E,
	0x5D, 0x36, 0x0D, 0x15, 0x38, 0x0F, 0x73, 0x2F, 0x35, 0x23, 0x25, 0x74,
	0x47, 0x09, 0x20, 0x08, 0x10, 0x2F, 0x17, 0x2D, 0x0C, 0x3A, 0x5F, 0x12,
	0x3D, 0x06, 0x6D, 0x26, 0x4E, 0x16, 0x01, 0x2D, 0x58, 0x59, 0x08, 0x06,
	0x73, 0x08, 0x18, 0x05, 0x3F, 0x0E, 0x2B, 0x08, 0x41, 0x25, 0x1A, 0x5F,
	0x58, 0x3C, 0x0E, 0x26, 0x3C, 0x36, 0x37, 0x5A, 0x7A, 0x47, 0x07, 0x1D,
	0x44, 0x71, 0x20, 0x31, 0x41, 0x40, 0x15, 0x47, 0x4E, 0x03, 0x39, 0x17,
	0x2A, 0x13, 0x14, 0x33, 0x05, 0x54, 0x10, 0x0B, 0x38, 0x01, 0x14, 0x2E,
	0x5F, 0x3D, 0x3A, 0x3F, 0x14, 0x5F, 0x25, 0x2C, 0x5A, 0x51, 0x5A, 0x25,
	0x0F, 0x19, 0x0F, 0x5E, 0x12, 0x74, 0x04, 0x4E, 0x41, 0x5B, 0x33, 0x5F,
	0x23, 0x22, 0x5F, 0x0D, 0x29, 0x18, 0x01, 0x31, 0x0C, 0x0A, 0x50, 0x1B,
	0x05, 0x03, 0x21, 0x51, 0x5A, 0x39, 0x38, 0x2D, 0x3B, 0x0A, 0x58, 0x2C,
	0x16, 0x17, 0x57, 0x20, 0x7B, 0x28, 0x00, 0x06, 0x02, 0x33, 0x2B, 0x55,
	0x1C, 0x13, 0x15, 0x1C, 0x4A, 0x08, 0x0F, 0x0A, 0x0F, 0x31, 0x05, 0x3C,
	0x12, 0x09, 0x18, 0x3F, 0x31, 0x7A, 0x2A, 0x0A, 0x17, 0x0F, 0x2D, 0x1E,
	0x04, 0x3A, 0x0D, 0x34, 0x1D, 0x0E, 0x0B, 0x2C, 0x25, 0x18, 0x29, 0x2A,
	0x38, 0x0A, 0x19, 0x27, 0x58, 0x23, 0x76, 0x02, 0x22, 0x0F, 0x08, 0x0A,
	0x5F, 0x12, 0x5E, 0x0D, 0x72, 0x3D, 0x12, 0x3B, 0x5F, 0x28, 0x01, 0x15,
	0x21, 0x23, 0x34, 0x5C, 0x23, 0x09, 0x33, 0x08, 0x23, 0x53, 0x39, 0x5C,
	0x2D, 0x0A, 0x19, 0x59, 0x05, 0x01, 0x05, 0x59, 0x04, 0x52, 0x73, 0x35,
	0x59, 0x01, 0x09, 0x75, 0x34, 0x29, 0x24, 0x3F, 0x12, 0x3E, 0x03, 0x37,
	0x07, 0x26, 0x43, 0x0A, 0x28, 0x06, 0x21, 0x2F, 0x0B, 0x5D, 0x39, 0x06,
	0x1D, 0x52, 0x0B, 0x0F, 0x2A, 0x28, 0x58, 0x17, 0x2E, 0x35, 0x2E, 0x55,
	0x5F, 0x20, 0x2E, 0x0F, 0x18, 0x25, 0x27, 0x15, 0x0A, 0x00, 0x59, 0x53,
	0x0A, 0x38, 0x06, 0x20, 0x59, 0x11, 0x18, 0x3B, 0x1A, 0x5B, 0x34, 0x09,
	0x39, 0x1A, 0x24, 0x06, 0x0B, 0x50, 0x14, 0x0E, 0x72, 0x55, 0x25, 0x3C,
	0x27, 0x2F, 0x0A, 0x2E, 0x37, 0x24, 0x69, 0x07, 0x04, 0x0F, 0x1B, 0x3A,
	0x23, 0x52, 0x5A, 0x25, 0x09, 0x26, 0x04, 0x0B, 0x21, 0x12, 0x58, 0x4E,
	0x28, 0x40, 0x26, 0x34, 0x11, 0x5B, 0x2F, 0x18, 0x2E, 0x56, 0x26, 0x24,
	0x0F, 0x5F, 0x0B, 0x19, 0x0C, 0x71, 0x2B, 0x26, 0x17, 0x59, 0x7B, 0x21,
	0x30, 0x0B, 0x5B, 0x70, 0x5C, 0x18, 0x5C, 0x04, 0x3B, 0x28, 0x24, 0x39,
	0x5C, 0x1A, 0x34, 0x51, 0x09, 0x27, 0x36, 0x22, 0x08, 0x56, 0x3F, 0x36,
	0x24, 0x00, 0x2D, 0x29, 0x2D, 0x0F, 0x36, 0x06, 0x00, 0x20, 0x24, 0x33,
	0x1F, 0x52, 0x07, 0x18, 0x29, 0x5F, 0x5E, 0x16, 0x36, 0x4E, 0x0B, 0x1D,
	0x1B, 0x5B, 0x1B, 0x05, 0x0F, 0x69, 0x08, 0x2E, 0x16, 0x1B, 0x76, 0x24,
	0x0F, 0x3F, 0x5F, 0x34, 0x1F, 0x11, 0x23, 0x08, 0x6D, 0x01, 0x34, 0x04,
	0x5A, 0x11, 0x1F, 0x14, 0x2B, 0x0C, 0x38, 0x5A, 0x0D, 0x3F, 0x03, 0x14,
	0x00, 0x35, 0x3D, 0x1F, 0x25, 0x28, 0x05, 0x28, 0x53, 0x2B, 0x2A, 0x19,
	0x21, 0x2C, 0x16, 0x19, 0x36, 0x3D, 0x12, 0x6D, 0x3D, 0x19, 0x19, 0x40,
	0x15, 0x2E, 0x1B, 0x1B, 0x1C, 0x70, 0x1D, 0x23, 0x00, 0x5B, 0x24, 0x0B,
	0x11, 0x17, 0x01, 0x18, 0x5B, 0x27, 0x0F, 0x26, 0x04, 0x5A, 0x28, 0x3E,
	0x39, 0x20, 0x1E, 0x0F, 0x1E, 0x5E, 0x16, 0x19, 0x0F, 0x23, 0x3F, 0x04,
	0x5A, 0x55, 0x2A, 0x2A, 0x16, 0x02, 0x09, 0x20, 0x25, 0x73, 0x25, 0x0F,
	0x3A, 0x58, 0x20, 0x26, 0x2E, 0x17, 0x3C, 0x77, 0x1E, 0x02, 0x04, 0x0A,
	0x14, 0x27, 0x06, 0x37, 0x00, 0x73, 0x16, 0x2A, 0x21, 0x40, 0x3A, 0x3F,
	0x13, 0x24, 0x32, 0x2E, 0x5E, 0x07, 0x2A, 0x28, 0x28, 0x39, 0x07, 0x3A,
	0x0C, 0x70, 0x58, 0x09, 0x3B, 0x28, 0x13, 0x5C, 0x30, 0x0A, 0x01, 0x11,
	0x35, 0x53, 0x5B, 0x5E, 0x29, 0x29, 0x12, 0x0B, 0x25, 0x0B, 0x28, 0x07,
	0x5E, 0x3F, 0x20, 0x28, 0x0F, 0x14, 0x05, 0x2F, 0x38, 0x0B, 0x22, 0x0F,
	0x0A, 0x2A, 0x55, 0x5B, 0x52, 0x1B, 0x0F, 0x4E, 0x58, 0x2F, 0x20, 0x25,
	0x26, 0x08, 0x5E, 0x18, 0x19, 0x04, 0x20, 0x13, 0x73, 0x1C, 0x54, 0x1A,
	0x13, 0x00, 0x58, 0x23, 0x18, 0x38, 0x33, 0x1A, 0x0F, 0x3A, 0x23, 0x69,
	0x19, 0x4A, 0x14, 0x32, 0x15, 0x2A, 0x34, 0x26, 0x2D, 0x00, 0x55, 0x56,
	0x29, 0x1C, 0x70, 0x02, 0x03, 0x5B, 0x26, 0x37, 0x19, 0x52, 0x02, 0x33,
	0x13, 0x2F, 0x33, 0x24, 0x33, 0x01, 0x04, 0x30, 0x58, 0x59, 0x7B, 0x43,
	0x38, 0x29, 0x2F, 0x30, 0x0E, 0x55, 0x1E, 0x25, 0x05, 0x18, 0x52, 0x5B,
	0x0E, 0x77, 0x0D, 0x0C, 0x19, 0x11, 0x38, 0x16, 0x20, 0x00, 0x59, 0x27,
	0x19, 0x05, 0x23, 0x3D, 0x75, 0x29, 0x19, 0x5C, 0x28, 0x71, 0x1A, 0x19,
	0x3C, 0x00, 0x0C, 0x14, 0x36, 0x1F, 0x3B, 0x70, 0x2F, 0x36, 0x3D, 0x19,
	0x25, 0x3A, 0x33, 0x2D, 0x24, 0x2C, 0x15, 0x1B, 0x08, 0x3A, 0x05, 0x1E,
	0x00, 0x37, 0x1F, 0x69, 0x07, 0x34, 0x08, 0x3D, 0x12, 0x2A, 0x13, 0x1B,
	0x3A, 0x70, 0x5C, 0x19, 0x1F, 0x23, 0x34, 0x14, 0x0A, 0x02, 0x04, 0x33,
	0x29, 0x15, 0x5E, 0x0F, 0x35, 0x34, 0x25, 0x29, 0x24, 0x16, 0x15, 0x32,
	0x3E, 0x3C, 0x2C, 0x0D, 0x34, 0x2A, 0x1B, 0x0C, 0x5E, 0x18, 0x04, 0x26,
	0x29, 0x54, 0x33, 0x28, 0x26, 0x0C, 0x5A, 0x58, 0x3F, 0x22, 0x35, 0x27,
	0x39, 0x56, 0x0F, 0x73, 0x2F, 0x50, 0x0A, 0x09, 0x08, 0x43, 0x26, 0x34,
	0x18, 0x07, 0x43, 0x2C, 0x3D, 0x1B, 0x23, 0x54, 0x35, 0x39, 0x31, 0x71,
	0x43, 0x13, 0x59, 0x12, 0x75, 0x16, 0x23, 0x1C, 0x58, 0x25, 0x22, 0x58,
	0x23, 0x21, 0x6D, 0x14, 0x05, 0x09, 0x03, 0x2B, 0x5D, 0x00, 0x1B, 0x5B,
	0x74, 0x3A, 0x58, 0x28, 0x53, 0x20, 0x3D, 0x4E, 0x05, 0x1B, 0x6D, 0x2B,
	0x36, 0x36, 0x03, 0x21, 0x2F, 0x0B, 0x20, 0x31, 0x21, 0x26, 0x0B, 0x0A,
	0x25, 0x28, 0x27, 0x04, 0x0D, 0x18, 0x33, 0x07, 0x2D, 0x57, 0x09, 0x3B,
	0x3C, 0x13, 0x26, 0x5D, 0x13, 0x38, 0x33, 0x0A, 0x0E, 0x11, 0x1E, 0x0C,
	0x1A, 0x52, 0x31, 0x18, 0x06, 0x56, 0x27, 0x30, 0x1B, 0x54, 0x34, 0x28,
	0x0A, 0x3A, 0x11, 0x2F, 0x0A, 0x3A, 0x3C, 0x27, 0x0C, 0x1B, 0x04, 0x0D,
	0x56, 0x29, 0x06, 0x31, 0x25, 0x29, 0x0F, 0x11, 0x6D, 0x06, 0x17, 0x0D,
	0x3A, 0x0E, 0x5E, 0x0B, 0x0A, 0x0E, 0x2E, 0x55, 0x03, 0x05, 0x3C, 0x3B,
	0x19, 0x4E, 0x21, 0x58, 0x76, 0x3B, 0x53, 0x3E, 0x07, 0x1B, 0x5C, 0x36,
	0x0D, 0x02, 0x13, 0x39, 0x39, 0x09, 0x2C, 0x26, 0x5A, 0x39, 0x29, 0x12,
	0x2E, 0x5D, 0x22, 0x0B, 0x2F, 0x69, 0x3C, 0x14, 0x58, 0x1D, 0x00, 0x2E,
	0x34, 0x1D, 0x1E, 0x09, 0x18, 0x25, 0x5B, 0x59, 0x70, 0x25, 0x56, 0x56,
	0x5C, 0x21, 0x1E, 0x51, 0x2F, 0x00, 0x0B, 0x06, 0x3B, 0x41, 0x3F, 0x13,
	0x00, 0x09, 0x36, 0x0F, 0x31, 0x39, 0x04, 0x18, 0x20, 0x32, 0x3E, 0x17,
	0x01, 0x3E, 0x16, 0x0E, 0x30, 0x38, 0x39, 0x1A, 0x08, 0x0C, 0x2A, 0x3F,
	0x2D, 0x3A, 0x12, 0x26, 0x1E, 0x17, 0x5F, 0x03, 0x3C, 0x38, 0x21, 0x3F,
	0x2B, 0x2B, 0x0C, 0x03, 0x09, 0x2D, 0x3D, 0x28, 0x1A, 0x39, 0x0C, 0x5F,
	0x2A, 0x38, 0x3C, 0x56, 0x2F, 0x53, 0x31, 0x35, 0x18, 0x58, 0x03, 0x31,
	0x22, 0x59, 0x0D, 0x12, 0x74, 0x0F, 0x38, 0x1C, 0x28, 0x0A, 0x0E, 0x33,
	0x08, 0x2D, 0x2B, 0x15, 0x27, 0x45, 0x3C, 0x71, 0x1F, 0x0C, 0x1D, 0x1B,
	0x0F, 0x35, 0x07, 0x22, 0x5D, 0x23, 0x0D, 0x10, 0x02, 0x09, 0x2A, 0x5B,
	0x2C, 0x56, 0x53, 0x2E, 0x20, 0x14, 0x1C, 0x29, 0x33, 0x18, 0x59, 0x2A,
	0x3A, 0x2F, 0x3B, 0x04, 0x1B, 0x23, 0x28, 0x3F, 0x2D, 0x5C, 0x23, 0x17,
	0x04, 0x2A, 0x1C, 0x44, 0x01, 0x1C, 0x57, 0x00, 0x44, 0x25, 0x1D, 0x04,
	0x01, 0x3C, 0x3A, 0x04, 0x0A, 0x3A, 0x32, 0x37, 0x28, 0x59, 0x2A, 0x44,
	0x0E, 0x0A, 0x22, 0x41, 0x08, 0x77, 0x5B, 0x55, 0x17, 0x3E, 0x04, 0x25,
	0x19, 0x3F, 0x5D, 0x6D, 0x20, 0x07, 0x2A, 0x44, 0x11, 0x1B, 0x06, 0x22,
	0x1C, 0x1A, 0x47, 0x28, 0x18, 0x1D, 0x06, 0x38, 0x04, 0x0B, 0x27, 0x7B,
	0x24, 0x54, 0x5A, 0x3E, 0x2E, 0x5A, 0x17, 0x14, 0x13, 0x09, 0x3B, 0x56,
	0x5E, 0x40, 0x03, 0x04, 0x20, 0x2F, 0x52, 0x75, 0x5C, 0x59, 0x3D, 0x18,
	0x69, 0x3D, 0x24, 0x16, 0x12, 0x3A, 0x58, 0x26, 0x1F, 0x02, 0x01, 0x55,
	0x24, 0x0C, 0x26, 0x7A, 0x25, 0x30, 0x04, 0x2A, 0x01, 0x5B, 0x07, 0x3C,
	0x2A, 0x26, 0x18, 0x1B, 0x2F, 0x3D, 0x2D, 0x0B, 0x58, 0x3B, 0x3A, 0x25,
	0x01, 0x53, 0x5B, 0x5E, 0x0C, 0x01, 0x06, 0x1F, 0x5E, 0x2D, 0x3F, 0x10,
	0x1E, 0x52, 0x08, 0x0B, 0x56, 0x1D, 0x0D, 0x18, 0x0F, 0x37, 0x28, 0x0F,
	0x15, 0x3F, 0x53, 0x2B, 0x12, 0x24, 0x5E, 0x13, 0x34, 0x1F, 0x23, 0x2F,
	0x18, 0x21, 0x21, 0x13, 0x36, 0x08, 0x04, 0x19, 0x72, 0x1D, 0x2F, 0x1B,
	0x31, 0x16, 0x0D, 0x34, 0x0D, 0x5C, 0x26, 0x09, 0x35, 0x1C, 0x0D, 0x2B,
	0x1D, 0x57, 0x2F, 0x0A, 0x23, 0x34, 0x34, 0x28, 0x52, 0x77, 0x18, 0x02,
	0x3F, 0x1B, 0x36, 0x19, 0x15, 0x45, 0x0E, 0x08, 0x39, 0x22, 0x38, 0x5E,
	0x03, 0x16, 0x20, 0x17, 0x0E, 0x21, 0x26, 0x14, 0x1A, 0x2D, 0x24, 0x38,
	0x28, 0x19, 0x5A, 0x0B, 0x1A, 0x17, 0x20, 0x2D, 0x30, 0x28, 0x3B, 0x24,
	0x05, 0x2F, 0x36, 0x19, 0x5B, 0x3C, 0x7B, 0x0E, 0x2E, 0x09, 0x5B, 0x74,
	0x2E, 0x57, 0x59, 0x2E, 0x29, 0x43, 0x04, 0x19, 0x39, 0x2F, 0x06, 0x29,
	0x58, 0x5F, 0x07, 0x55, 0x16, 0x1E, 0x28, 0x13, 0x2E, 0x38, 0x3B, 0x2E,
	0x36, 0x34, 0x52, 0x2F, 0x5C, 0x32, 0x0E, 0x15, 0x2F, 0x09, 0x35, 0x38,
	0x14, 0x3E, 0x1C, 0x03, 0x39, 0x27, 0x21, 0x28, 0x04, 0x09, 0x09, 0x0A,
	0x2D, 0x2A, 0x20, 0x24, 0x5A, 0x19, 0x29, 0x39, 0x37, 0x5F, 0x01, 0x0E,
	0x1B, 0x17, 0x16, 0x1E, 0x0D, 0x1F, 0x27, 0x58, 0x58, 0x04, 0x08, 0x32,
	0x3D, 0x13, 0x06, 0x00, 0x04, 0x56, 0x1C, 0x2D, 0x23, 0x22, 0x1E, 0x1A,
	0x73, 0x43, 0x32, 0x0B, 0x04, 0x35, 0x55, 0x50, 0x07, 0x59, 0x24, 0x5D,
	0x28, 0x39, 0x13, 0x69, 0x5D, 0x0E, 0x0B, 0x5B, 0x08, 0x5E, 0x08, 0x41,
	0x1F, 0x73, 0x3A, 0x56, 0x1A, 0x12, 0x69, 0x01, 0x16, 0x57, 0x39, 0x7A,
	0x3F, 0x24, 0x24, 0x0C, 0x12, 0x2D, 0x0C, 0x2C, 0x0D, 0x71, 0x3B, 0x35,
	0x18, 0x18, 0x28, 0x59, 0x14, 0x57, 0x0C, 0x2A, 0x5B, 0x55, 0x1F, 0x1B,
	0x0E, 0x3C, 0x05, 0x27, 0x21, 0x20, 0x18, 0x16, 0x2B, 0x0D, 0x18, 0x26,
	0x36, 0x04, 0x05, 0x7A, 0x0E, 0x08, 0x58, 0x0E, 0x70, 0x0F, 0x2E, 0x5F,
	0x44, 0x33, 0x1E, 0x05, 0x5C, 0x20, 0x07, 0x07, 0x07, 0x5D, 0x0A, 0x15,
	0x1C, 0x26, 0x3F, 0x58, 0x11, 0x1A, 0x54, 0x2C, 0x25, 0x0A, 0x06, 0x58,
	0x3F, 0x25, 0x08, 0x3F, 0x02, 0x23, 0x1F, 0x08, 0x5D, 0x00, 0x08, 0x20,
	0x10, 0x5B, 0x23, 0x22, 0x25, 0x72, 0x14, 0x33, 0x04, 0x2E, 0x13, 0x1D,
	0x32, 0x0D, 0x11, 0x3A, 0x3E, 0x38, 0x5C, 0x1E, 0x37, 0x34, 0x33, 0x45,
	0x2E, 0x10, 0x1F, 0x4E, 0x3D, 0x58, 0x0B, 0x09, 0x20, 0x2D, 0x1B, 0x2F,
	0x5A, 0x53, 0x19, 0x25, 0x11, 0x08, 0x22, 0x2C, 0x3D, 0x31, 0x2B, 0x38,
	0x08, 0x18, 0x11, 0x06, 0x0C, 0x59, 0x20, 0x28, 0x1F, 0x16, 0x2A, 0x5A,
	0x6D, 0x3C, 0x14, 0x09, 0x20, 0x01, 0x39, 0x54, 0x5E, 0x0C, 0x06, 0x2F,
	0x52, 0x0F, 0x27, 0x71, 0x0E, 0x50, 0x3F, 0x3B, 0x03, 0x0D, 0x10, 0x1C,
	0x40, 0x00, 0x03, 0x39, 0x18, 0x3C, 0x3A, 0x2F, 0x08, 0x08, 0x33, 0x2D,
	0x2F, 0x23, 0x29, 0x1D, 0x33, 0x1C, 0x37, 0x25, 0x06, 0x29, 0x2B, 0x59,
	0x41, 0x39, 0x34, 0x02, 0x27, 0x1D, 0x2D, 0x34, 0x06, 0x35, 0x06, 0x5D,
	0x25, 0x27, 0x2D, 0x18, 0x52, 0x0C, 0x47, 0x05, 0x20, 0x2D, 0x0B, 0x47,
	0x0E, 0x0F, 0x5D, 0x69, 0x03, 0x27, 0x41, 0x39, 0x13, 0x0D, 0x07, 0x19,
	0x5D, 0x06, 0x08, 0x2C, 0x14, 0x2F, 0x09, 0x25, 0x36, 0x0D, 0x5C, 0x08,
	0x29, 0x37, 0x2C, 0x01, 0x32, 0x1F, 0x54, 0x02, 0x1B, 0x77, 0x2E, 0x4E,
	0x5A, 0x3D, 0x18, 0x3B, 0x25, 0x38, 0x39, 0x73, 0x0A, 0x13, 0x03, 0x28,
	0x0B, 0x02, 0x3B, 0x21, 0x05, 0x33, 0x0A, 0x03, 0x58, 0x5A, 0x75, 0x06,
	0x38, 0x3B, 0x0F, 0x20, 0x54, 0x20, 0x3D, 0x3B, 0x27, 0x0B, 0x59, 0x01,
	0x01, 0x2E, 0x20, 0x0D, 0x0F, 0x0A, 0x3A, 0x25, 0x02, 0x34, 0x3C, 0x06,
	0x18, 0x2A, 0x5E, 0x52, 0x7A, 0x20, 0x36, 0x3E, 0x5D, 0x0E, 0x35, 0x33,
	0x5C, 0x0C, 0x74, 0x35, 0x54, 0x14, 0x0F, 0x7B, 0x0F, 0x09, 0x20, 0x3C,
	0x06, 0x5B, 0x0E, 0x37, 0x1E, 0x15, 0x39, 0x52, 0x00, 0x0E, 0x08, 0x03,
	0x06, 0x01, 0x2A, 0x04, 0x0B, 0x00, 0x5E, 0x58, 0x0A, 0x18, 0x55, 0x17,
	0x0F, 0x26, 0x05, 0x50, 0x0C, 0x1C, 0x76, 0x38, 0x37, 0x45, 0x2C, 0x32,
	0x29, 0x00, 0x00, 0x12, 0x07, 0x29, 0x56, 0x06, 0x0C, 0x0E, 0x54, 0x08,
	0x41, 0x39, 0x15, 0x1C, 0x1B, 0x0C, 0x04, 0x24, 0x14, 0x55, 0x27, 0x5A,
	0x0C, 0x5B, 0x26, 0x2A, 0x1F, 0x2C, 0x18, 0x19, 0x39, 0x33, 0x28, 0x43,
	0x50, 0x41, 0x2F, 0x2C, 0x21, 0x24, 0x06, 0x0D, 0x37, 0x0B, 0x2C, 0x58,
	0x09, 0x29, 0x09, 0x54, 0x3C, 0x5E, 0x14, 0x19, 0x11, 0x0F, 0x52, 0x70,
	0x27, 0x0F, 0x59, 0x3F, 0x71, 0x26, 0x17, 0x37, 0x5F, 0x25, 0x1D, 0x00,
	0x2B, 0x20, 0x32, 0x5D, 0x24, 0x2B, 0x2C, 0x75, 0x09, 0x00, 0x2A, 0x29,
	0x34, 0x09, 0x56, 0x59, 0x5E, 0x16, 0x47, 0x4E, 0x37, 0x19, 0x77, 0x0A,
	0x2C, 0x1F, 0x2A, 0x36, 0x5C, 0x06, 0x3B, 0x3F, 0x70, 0x3F, 0x05, 0x02,
	0x5B, 0x0A, 0x3A, 0x59, 0x23, 0x0D, 0x31, 0x27, 0x51, 0x17, 0x2C, 0x06,
	0x3F, 0x37, 0x41, 0x08, 0x0C, 0x3A, 0x2C, 0x1B, 0x12, 0x2F, 0x0D, 0x11,
	0x07, 0x40, 0x0A, 0x06, 0x00, 0x1B, 0x2E, 0x1B, 0x5C, 0x11, 0x3D, 0x23,
	0x71, 0x3D, 0x2D, 0x3E, 0x33, 0x71, 0x59, 0x28, 0x2C, 0x1D, 0x1B, 0x01,
	0x58, 0x34, 0x32, 0x04, 0x5A, 0x29, 0x18, 0x06, 0x6D, 0x26, 0x17, 0x27,
	0x5A, 0x21, 0x0D, 0x16, 0x28, 0x1F, 0x12, 0x1E, 0x23, 0x00, 0x5B, 0x27,
	0x1B, 0x2B, 0x24, 0x2E, 0x12, 0x15, 0x4A, 0x20, 0x25, 0x7B, 0x20, 0x53,
	0x58, 0x1C, 0x0A, 0x5D, 0x20, 0x1D, 0x03, 0x15, 0x59, 0x4A, 0x08, 0x5D,
	0x26, 0x55, 0x30, 0x41, 0x23, 0x25, 0x38, 0x51, 0x17, 0x01, 0x38, 0x23,
	0x31, 0x56, 0x5A, 0x29, 0x1D, 0x36, 0x3C, 0x0A, 0x36, 0x05, 0x35, 0x18,
	0x3E, 0x28, 0x14, 0x22, 0x1D, 0x11, 0x12, 0x5F, 0x32, 0x07, 0x01, 0x2F,
	0x14, 0x4E, 0x5A, 0x5C, 0x2A, 0x47, 0x07, 0x18, 0x2D, 0x26, 0x0A, 0x06,
	0x04, 0x01, 0x0D, 0x09, 0x36, 0x26, 0x05, 0x0A, 0x3D, 0x2E, 0x1D, 0x39,
	0x35, 0x1E, 0x56, 0x56, 0x1D, 0x1B, 0x43, 0x52, 0x3D, 0x02, 0x14, 0x28,
	0x11, 0x24, 0x22, 0x2F, 0x3F, 0x39, 0x17, 0x01, 0x14, 0x0E, 0x52, 0x06,
	0x25, 0x2F, 0x38, 0x04, 0x39, 0x5D, 0x29, 0x02, 0x37, 0x0C, 0x0E, 0x1A,
	0x28, 0x39, 0x21, 0x33, 0x38, 0x21, 0x08, 0x39, 0x38, 0x2E, 0x20, 0x02,
	0x5A, 0x03, 0x31, 0x2E, 0x58, 0x0F, 0x2E, 0x09, 0x14, 0x06, 0x14, 0x12,
	0x28, 0x3B, 0x0A, 0x3D, 0x29, 0x0E, 0x0A, 0x2C, 0x27, 0x24, 0x07, 0x19,
	0x52, 0x14, 0x05, 0x21, 0x34, 0x3B, 0x25, 0x28, 0x71, 0x06, 0x10, 0x1B,
	0x0F, 0x03, 0x2B, 0x37, 0x24, 0x2A, 0x16, 0x3A, 0x26, 0x5A, 0x23, 0x13,
	0x28, 0x4E, 0x26, 0x53, 0x2B, 0x55, 0x2A, 0x0D, 0x02, 0x2E, 0x5D, 0x16,
	0x17, 0x01, 0x0D, 0x15, 0x12, 0x37, 0x32, 0x27, 0x0F, 0x3B, 0x39, 0x3A,
	0x7B, 0x1A, 0x1B, 0x23, 0x27, 0x73, 0x29, 0x28, 0x59, 0x5D, 0x18, 0x1E,
	0x2F, 0x37, 0x27, 0x33, 0x0D, 0x22, 0x3D, 0x40, 0x0C, 0x3A, 0x12, 0x1E,
	0x01, 0x04, 0x0D, 0x52, 0x22, 0x5B, 0x7B, 0x18, 0x0C, 0x34, 0x23, 0x0C,
	0x5E, 0x08, 0x3B, 0x3D, 0x73, 0x2F, 0x03, 0x5B, 0x1B, 0x30, 0x3F, 0x36,
	0x03, 0x39, 0x2E, 0x5A, 0x33, 0x3B, 0x11, 0x15, 0x02, 0x05, 0x5B, 0x3A,
	0x37, 0x0F, 0x0C, 0x16, 0x1D, 0x75, 0x0F, 0x52, 0x3D, 0x3D, 0x3A, 0x06,
	0x09, 0x19, 0x09, 0x01, 0x39, 0x0E, 0x06, 0x3B, 0x2D, 0x03, 0x2C, 0x3B,
	0x27, 0x11, 0x47, 0x10, 0x5C, 0x58, 0x6D, 0x0F, 0x0C, 0x25, 0x09, 0x26,
	0x29, 0x55, 0x5C, 0x58, 0x0F, 0x47, 0x17, 0x06, 0x02, 0x70, 0x36, 0x25,
	0x5F, 0x58, 0x30, 0x1D, 0x33, 0x56, 0x52, 0x12, 0x3A, 0x23, 0x5B, 0x2C,
	0x2C, 0x14, 0x0B, 0x14, 0x13, 0x0D, 0x3B, 0x15, 0x05, 0x1D, 0x3B, 0x3E,
	0x30, 0x19, 0x5C, 0x09, 0x20, 0x39, 0x25, 0x01, 0x0B, 0x5A, 0x08, 0x0A,
	0x23, 0x38, 0x14, 0x53, 0x23, 0x38, 0x2B, 0x1D, 0x51, 0x0D, 0x08, 0x0C,
	0x2E, 0x04, 0x22, 0x2C, 0x0C, 0x07, 0x05, 0x02, 0x27, 0x76, 0x58, 0x54,
	0x37, 0x1F, 0x17, 0x5E, 0x31, 0x3E, 0x05, 0x14, 0x59, 0x0A, 0x16, 0x1D,
	0x07, 0x5A, 0x15, 0x39, 0x1C, 0x2F, 0x23, 0x23, 0x23, 0x1A, 0x24, 0x3F,
	0x55, 0x3A, 0x5A, 0x7B, 0x1A, 0x13, 0x06, 0x1A, 0x0C, 0x47, 0x13, 0x38,
	0x5E, 0x74, 0x3C, 0x18, 0x0C, 0x0F, 0x71, 0x06, 0x0A, 0x26, 0x08, 0x74,
	0x27, 0x0F, 0x0D, 0x32, 0x1B, 0x2F, 0x2D, 0x03, 0x07, 0x12, 0x0A, 0x15,
	0x59, 0x23, 0x16, 0x25, 0x39, 0x14, 0x07, 0x70, 0x0A, 0x0D, 0x1B, 0x3A,
	0x24, 0x5D, 0x10, 0x1D, 0x1D, 0x2F, 0x1D, 0x30, 0x19, 0x09, 0x01, 0x0B,
	0x22, 0x3A, 0x5B, 0x30, 0x18, 0x2D, 0x38, 0x24, 0x24, 0x09, 0x57, 0x5B,
	0x5E, 0x3B, 0x58, 0x30, 0x38, 0x5A, 0x70, 0x0E, 0x10, 0x0F, 0x53, 0x03,
	0x23, 0x1B, 0x34, 0x03, 0x0D, 0x22, 0x52, 0x3A, 0x1E, 0x31, 0x54, 0x09,
	0x1A, 0x5D, 0x07, 0x20, 0x2F, 0x26, 0x00, 0x12, 0x3A, 0x2E, 0x5B, 0x0E,
	0x09, 0x08, 0x06, 0x5B, 0x0F, 0x29, 0x2F, 0x0A, 0x2C, 0x5C, 0x7B, 0x5C,
	0x55, 0x1E, 0x5D, 0x38, 0x3D, 0x54, 0x05, 0x1D, 0x3B, 0x20, 0x12, 0x1C,
	0x0E, 0x72, 0x05, 0x19, 0x36, 0x11, 0x17, 0x21, 0x3B, 0x37, 0x28, 0x71,
	0x19, 0x51, 0x3C, 0x08, 0x7B, 0x3B, 0x24, 0x1F, 0x3B, 0x23, 0x3B, 0x2D,
	0x1F, 0x5D, 0x76, 0x0A, 0x25, 0x24, 0x05, 0x01, 0x07, 0x34, 0x28, 0x0F,
	0x7A, 0x2F, 0x15, 0x0F, 0x5E, 0x30, 0x2A, 0x39, 0x09, 0x0E, 0x32, 0x5D,
	0x39, 0x3F, 0x31, 0x0C, 0x2B, 0x58, 0x5B, 0x23, 0x20, 0x3B, 0x2C, 0x3A,
	0x40, 0x2E, 0x2A, 0x18, 0x20, 0x20, 0x16, 0x3D, 0x58, 0x45, 0x00, 0x34,
	0x19, 0x0A, 0x27, 0x5A, 0x2D, 0x22, 0x15, 0x5B, 0x58, 0x16, 0x5C, 0x53,
	0x5F, 0x24, 0x37, 0x5C, 0x3B, 0x1B, 0x26, 0x04, 0x3A, 0x1B, 0x2A, 0x00,
	0x29, 0x28, 0x58, 0x5D, 0x00, 0x05, 0x09, 0x28, 0x27, 0x1D, 0x05, 0x22,
	0x03, 0x5F, 0x11, 0x00, 0x1B, 0x53, 0x20, 0x05, 0x09, 0x1E, 0x0F, 0x1C,
	0x28, 0x76, 0x3F, 0x17, 0x00, 0x0F, 0x1B, 0x28, 0x52, 0x07, 0x0A, 0x20,
	0x0E, 0x18, 0x5B, 0x1C, 0x69, 0x3D, 0x30, 0x2C, 0x0F, 0x75, 0x58, 0x0D,
	0x37, 0x0D, 0x31, 0x5B, 0x0D, 0x5C, 0x26, 0x07, 0x03, 0x02, 0x05, 0x1B,
	0x75, 0x58, 0x00, 0x06, 0x40, 0x37, 0x2A, 0x2C, 0x39, 0x04, 0x32, 0x59,
	0x3B, 0x17, 0x27, 0x14, 0x5C, 0x04, 0x59, 0x06, 0x03, 0x1F, 0x2C, 0x57,
	0x01, 0x2C, 0x0F, 0x16, 0x24, 0x0F, 0x7A, 0x25, 0x14, 0x3C, 0x2C, 0x09,
	0x19, 0x33, 0x23, 0x3E, 0x33, 0x0E, 0x27, 0x21, 0x31, 0x1B, 0x59, 0x2F,
	0x17, 0x3D, 0x76, 0x1E, 0x15, 0x2A, 0x1F, 0x7B, 0x25, 0x4E, 0x21, 0x1F,
	0x0B, 0x3B, 0x4E, 0x2F, 0x25, 0x31, 0x5D, 0x0F, 0x28, 0x24, 0x06, 0x5B,
	0x57, 0x0D, 0x13, 0x36, 0x14, 0x29, 0x5E, 0x0C, 0x20, 0x00, 0x11, 0x03,
	0x26, 0x0D, 0x0D, 0x30, 0x06, 0x11, 0x28, 0x00, 0x36, 0x57, 0x26, 0x74,
	0x20, 0x07, 0x20, 0x1A, 0x33, 0x2A, 0x30, 0x41, 0x1B, 0x74, 0x1F, 0x09,
	0x3A, 0x3C, 0x21, 0x5E, 0x28, 0x0C, 0x1E, 0x2F, 0x1B, 0x2F, 0x3A, 0x40,
	0x2C, 0x47, 0x4E, 0x09, 0x5B, 0x35, 0x15, 0x59, 0x2F, 0x0C, 0x7A, 0x55,
	0x12, 0x09, 0x03, 0x2C, 0x09, 0x36, 0x3D, 0x03, 0x0D, 0x5C, 0x24, 0x1A,
	0x27, 0x0C, 0x1D, 0x03, 0x28, 0x2A, 0x72, 0x3C, 0x59, 0x0C, 0x52, 0x0B,
	0x5C, 0x33, 0x16, 0x1B, 0x2C, 0x3F, 0x52, 0x16, 0x44, 0x29, 0x34, 0x2D,
	0x17, 0x58, 0x2A, 0x2A, 0x0F, 0x1F, 0x25, 0x3B, 0x3C, 0x4A, 0x5B, 0x2C,
	0x35, 0x5F, 0x09, 0x06, 0x1D, 0x35, 0x20, 0x2D, 0x57, 0x1E, 0x74, 0x5D,
	0x4A, 0x3E, 0x0D, 0x7B, 0x2E, 0x00, 0x3F, 0x2F, 0x30, 0x1B, 0x15, 0x39,
	0x1F, 0x69, 0x22, 0x28, 0x5E, 0x04, 0x76, 0x21, 0x4A, 0x27, 0x0E, 0x25,
	0x22, 0x18, 0x19, 0x2A, 0x15, 0x03, 0x0B, 0x18, 0x3E, 0x08, 0x3A, 0x36,
	0x04, 0x2C, 0x2A, 0x0B, 0x38, 0x26, 0x28, 0x29, 0x0E, 0x50, 0x21, 0x00,
	0x08, 0x2D, 0x08, 0x37, 0x2A, 0x05, 0x15, 0x50, 0x2A, 0x0A, 0x2D, 0x2A,
	0x26, 0x00, 0x20, 0x3B, 0x5C, 0x58, 0x01, 0x1A, 0x2D, 0x5F, 0x55, 0x0F,
	0x00, 0x12, 0x15, 0x0B, 0x16, 0x03, 0x24, 0x05, 0x06, 0x09, 0x3F, 0x27,
	0x18, 0x37, 0x39, 0x38, 0x2F, 0x3A, 0x53, 0x27, 0x18, 0x34, 0x2F, 0x2E,
	0x36, 0x22, 0x7B, 0x43, 0x50, 0x2D, 0x03, 0x76, 0x04, 0x2A, 0x08, 0x5E,
	0x38, 0x1A, 0x18, 0x3A, 0x5F, 0x32, 0x1C, 0x23, 0x19, 0x2F, 0x08, 0x3A,
	0x28, 0x22, 0x28, 0x11, 0x21, 0x0F, 0x29, 0x18, 0x21, 0x23, 0x2B, 0x0A,
	0x0F, 0x27, 0x5B, 0x02, 0x5C, 0x0E, 0x6D, 0x35, 0x12, 0x39, 0x32, 0x2A,
	0x5A, 0x06, 0x3D, 0x05, 0x36, 0x3E, 0x2E, 0x58, 0x0F, 0x10, 0x28, 0x37,
	0x0B, 0x3A, 0x7B, 0x29, 0x02, 0x06, 0x0E, 0x2A, 0x0A, 0x57, 0x0D, 0x21,
	0x03, 0x1F, 0x55, 0x24, 0x02, 0x36, 0x5F, 0x18, 0x0D, 0x3D, 0x2E, 0x5D,
	0x18, 0x37, 0x0F, 0x26, 0x21, 0x15, 0x59, 0x5F, 0x1B, 0x21, 0x29, 0x1B,
	0x2F, 0x72, 0x5F, 0x54, 0x2D, 0x0D, 0x38, 0x43, 0x34, 0x09, 0x1B, 0x33,
	0x2A, 0x11, 0x0B, 0x1C, 0x0A, 0x08, 0x53, 0x57, 0x23, 0x75, 0x27, 0x55,
	0x0A, 0x05, 0x1B, 0x58, 0x3B, 0x0D, 0x59, 0x73, 0x1F, 0x52, 0x21, 0x5D,
	0x0F, 0x02, 0x2A, 0x2B, 0x5B, 0x71, 0x54, 0x29, 0x14, 0x01, 0x6D, 0x5F,
	0x27, 0x23, 0x23, 0x21, 0x3E, 0x38, 0x56, 0x2A, 0x31, 0x19, 0x24, 0x22,
	0x3B, 0x1B, 0x27, 0x55, 0x5E, 0x31, 0x71, 0x1E, 0x29, 0x06, 0x2F, 0x2C,
	0x2E, 0x08, 0x3B, 0x2F, 0x76, 0x1F, 0x1B, 0x25, 0x1D, 0x10, 0x03, 0x1B,
	0x20, 0x03, 0x29, 0x0D, 0x15, 0x16, 0x2E, 0x36, 0x23, 0x0E, 0x09, 0x24,
	0x76, 0x02, 0x3B, 0x2F, 0x58, 0x07, 0x55, 0x09, 0x24, 0x06, 0x18, 0x14,
	0x22, 0x45, 0x03, 0x38, 0x16, 0x08, 0x22, 0x1F, 0x06, 0x2A, 0x2E, 0x5E,
	0x3A, 0x70, 0x58, 0x09, 0x16, 0x2F, 0x33, 0x2E, 0x30, 0x5C, 0x5D, 0x11,
	0x2D, 0x19, 0x09, 0x25, 0x1A, 0x03, 0x4A, 0x02, 0x2F, 0x13, 0x3E, 0x17,
	0x25, 0x1B, 0x74, 0x25, 0x19, 0x2A, 0x3A, 0x2E, 0x5F, 0x2B, 0x2A, 0x3B,
	0x21, 0x1A, 0x0E, 0x08, 0x11, 0x18, 0x5D, 0x02, 0x05, 0x27, 0x24, 0x22,
	0x55, 0x3A, 0x5B, 0x05, 0x07, 0x14, 0x0C, 0x39, 0x1A, 0x2E, 0x14, 0x01,
	0x18, 0x10, 0x58, 0x57, 0x0A, 0x53, 0x11, 0x54, 0x2C, 0x07, 0x28, 0x2E,
	0x16, 0x07, 0x29, 0x0E, 0x38, 0x1D, 0x0C, 0x59, 0x33, 0x0F, 0x04, 0x03,
	0x0B, 0x24, 0x75, 0x54, 0x50, 0x5A, 0x25, 0x32, 0x1A, 0x16, 0x18, 0x25,
	0x20, 0x27, 0x26, 0x08, 0x03, 0x13, 0x1D, 0x10, 0x1A, 0x1B, 0x1A, 0x00,
	0x27, 0x2D, 0x11, 0x1B, 0x3E, 0x19, 0x57, 0x1F, 0x70, 0x47, 0x26, 0x01,
	0x3B, 0x0B, 0x5F, 0x58, 0x17, 0x12, 0x07, 0x47, 0x29, 0x0F, 0x11, 0x23,
	0x26, 0x14, 0x45, 0x3D, 0x7B, 0x14, 0x35, 0x27, 0x5C, 0x1A, 0x36, 0x19,
	0x5D, 0x3D, 0x20, 0x25, 0x18, 0x07, 0x5F, 0x0A, 0x09, 0x14, 0x58, 0x23,
	0x1A, 0x47, 0x07, 0x01, 0x09, 0x3A, 0x16, 0x18, 0x37, 0x08, 0x23, 0x1F,
	0x28, 0x57, 0x0D, 0x09, 0x23, 0x4E, 0x26, 0x28, 0x29, 0x07, 0x2F, 0x04,
	0x00, 0x23, 0x26, 0x20, 0x5C, 0x2E, 0x27, 0x08, 0x17, 0x5A, 0x07, 0x27,
	0x59, 0x13, 0x0D, 0x1D, 0x27, 0x3E, 0x26, 0x3A, 0x1D, 0x70, 0x22, 0x23,
	0x07, 0x27, 0x30, 0x19, 0x58, 0x1D, 0x1B, 0x27, 0x38, 0x31, 0x1D, 0x03,
	0x26, 0x5F, 0x59, 0x41, 0x1B, 0x70, 0x54, 0x24, 0x5B, 0x2F, 0x71, 0x5A,
	0x2B, 0x57, 0x19, 0x3A, 0x29, 0x50, 0x04, 0x1A, 0x6D, 0x07, 0x58, 0x09,
	0x40, 0x26, 0x00, 0x0F, 0x39, 0x28, 0x30, 0x1F, 0x24, 0x59, 0x2C, 0x72,
	0x24, 0x0F, 0x14, 0x3B, 0x09, 0x3F, 0x1B, 0x23, 0x23, 0x14, 0x43, 0x33,
	0x37, 0x13, 0x09, 0x1E, 0x07, 0x19, 0x05, 0x26, 0x5F, 0x27, 0x5B, 0x5A,
	0x10, 0x27, 0x16, 0x1F, 0x03, 0x0B, 0x08, 0x35, 0x3A, 0x3E, 0x0E, 0x59,
	0x22, 0x22, 0x38, 0x16, 0x20, 0x34, 0x45, 0x02, 0x0D, 0x14, 0x4A, 0x28,
	0x18, 0x2D, 0x14, 0x35, 0x14, 0x07, 0x35, 0x3C, 0x57, 0x3E, 0x53, 0x35,
	0x39, 0x35, 0x0C, 0x3E, 0x27, 0x26, 0x14, 0x2B, 0x2A, 0x27, 0x08, 0x0B,
	0x09, 0x0D, 0x6D, 0x0A, 0x07, 0x14, 0x1D, 0x15, 0x0E, 0x05, 0x58, 0x04,
	0x18, 0x55, 0x50, 0x29, 0x59, 0x3A, 0x27, 0x52, 0x26, 0x53, 0x12, 0x47,
	0x37, 0x08, 0x3E, 0x30, 0x5D, 0x0D, 0x28, 0x3C, 0x34, 0x14, 0x52, 0x1C,
	0x20, 0x0F, 0x1A, 0x13, 0x39, 0x3E, 0x24, 0x3E, 0x4E, 0x09, 0x02, 0x07,
	0x25, 0x2A, 0x41, 0x28, 0x13, 0x03, 0x26, 0x56, 0x1A, 0x71, 0x25, 0x03,
	0x07, 0x01, 0x73, 0x07, 0x04, 0x29, 0x03, 0x3A, 0x38, 0x52, 0x2C, 0x44,
	0x29, 0x18, 0x54, 0x02, 0x2D, 0x07, 0x0F, 0x32, 0x58, 0x12, 0x07, 0x3D,
	0x31, 0x2F, 0x2D, 0x1A, 0x21, 0x59, 0x3F, 0x44, 0x00, 0x2E, 0x1B, 0x1E,
	0x3A, 0x20, 0x07, 0x37, 0x1B, 0x1C, 0x0A, 0x1B, 0x31, 0x41, 0x32, 0x07,
	0x5A, 0x20, 0x25, 0x24, 0x3B, 0x1D, 0x2F, 0x05, 0x5A, 0x69, 0x0F, 0x03,
	0x06, 0x40, 0x70, 0x5C, 0x38, 0x24, 0x0D, 0x28, 0x0D, 0x15, 0x1E, 0x28,
	0x0D, 0x28, 0x0A, 0x04, 0x02, 0x21, 0x14, 0x12, 0x59, 0x3B, 0x75, 0x21,
	0x56, 0x45, 0x2F, 0x10, 0x29, 0x35, 0x19, 0x5B, 0x73, 0x20, 0x26, 0x09,
	0x53, 0x23, 0x0D, 0x0F, 0x06, 0x1A, 0x09, 0x24, 0x23, 0x3D, 0x0D, 0x0D,
	0x35, 0x2B, 0x14, 0x3C, 0x07, 0x43, 0x23, 0x45, 0x0D, 0x2E, 0x2D, 0x05,
	0x5B, 0x07, 0x13, 0x3B, 0x0C, 0x1F, 0x40, 0x14, 0x3F, 0x0A, 0x16, 0x1D,
	0x0B, 0x5E, 0x29, 0x45, 0x0F, 0x2E, 0x2A, 0x54, 0x0F, 0x03, 0x00, 0x0E,
	0x55, 0x37, 0x09, 0x72, 0x36, 0x1B, 0x18, 0x07, 0x07, 0x28, 0x25, 0x29,
	0x03, 0x04, 0x06, 0x17, 0x1D, 0x2F, 0x34, 0x09, 0x19, 0x5E, 0x5C, 0x28,
	0x07, 0x15, 0x1D, 0x20, 0x30, 0x21, 0x04, 0x3F, 0x01, 0x26, 0x14, 0x14,
	0x41, 0x5B, 0x28, 0x03, 0x2B, 0x5C, 0x5A, 0x0D, 0x1A, 0x2C, 0x04, 0x5A,
	0x21, 0x5B, 0x04, 0x56, 0x2F, 0x6D, 0x1F, 0x28, 0x1D, 0x2C, 0x31, 0x1E,
	0x2F, 0x23, 0x18, 0x0A, 0x29, 0x26, 0x1B, 0x1D, 0x2B, 0x5D, 0x09, 0x45,
	0x06, 0x73, 0x3C, 0x14, 0x01, 0x0A, 0x27, 0x08, 0x4A, 0x5A, 0x2D, 0x38,
	0x1C, 0x3B, 0x5C, 0x0F, 0x16, 0x01, 0x26, 0x26, 0x2E, 0x3B, 0x0A, 0x31,
	0x0C, 0x1D, 0x2E, 0x28, 0x17, 0x27, 0x52, 0x1B, 0x0A, 0x24, 0x21, 0x07,
	0x01, 0x21, 0x24, 0x04, 0x2D, 0x29, 0x02, 0x55, 0x2B, 0x22, 0x28, 0x1C,
	0x00, 0x0B, 0x08, 0x71, 0x54, 0x20, 0x59, 0x28, 0x26, 0x5B, 0x0B, 0x05,
	0x01, 0x76, 0x02, 0x09, 0x04, 0x5C, 0x05, 0x09, 0x28, 0x16, 0x11, 0x38,
	0x20, 0x59, 0x17, 0x52, 0x2F, 0x1E, 0x06, 0x37, 0x32, 0x2F, 0x5A, 0x27,
	0x14, 0x58, 0x71, 0x28, 0x04, 0x06, 0x0D, 0x1A, 0x3D, 0x54, 0x04, 0x0C,
	0x2A, 0x09, 0x56, 0x02, 0x2D, 0x2C, 0x0E, 0x29, 0x0B, 0x18, 0x2A, 0x3B,
	0x50, 0x05, 0x25, 0x03, 0x07, 0x2E, 0x26, 0x5F, 0x14, 0x27, 0x25, 0x0D,
	0x28, 0x6D, 0x3C, 0x58, 0x03, 0x2C, 0x2A, 0x5E, 0x0E, 0x06, 0x5A, 0x72,
	0x05, 0x30, 0x05, 0x5E, 0x2D, 0x28, 0x05, 0x0A, 0x33, 0x00, 0x00, 0x26,
	0x18, 0x3A, 0x10, 0x5B, 0x33, 0x3F, 0x26, 0x2E, 0x25, 0x56, 0x58, 0x29,
	0x73, 0x1B, 0x4A, 0x23, 0x11, 0x13, 0x54, 0x15, 0x1A, 0x39, 0x24, 0x07,
	0x15, 0x38, 0x26, 0x75, 0x2D, 0x18, 0x45, 0x59, 0x35, 0x55, 0x06, 0x2A,
	0x22, 0x35, 0x47, 0x4A, 0x1E, 0x3E, 0x17, 0x21, 0x29, 0x27, 0x28, 0x01,
	0x54, 0x29, 0x57, 0x3B, 0x28, 0x2E, 0x15, 0x16, 0x26, 0x0F, 0x03, 0x31,
	0x22, 0x0D, 0x2C, 0x29, 0x2A, 0x3B, 0x28, 0x36, 0x27, 0x59, 0x37, 0x44,
	0x01, 0x0B, 0x27, 0x1C, 0x5B, 0x08, 0x2B, 0x4E, 0x3A, 0x5A, 0x35, 0x34,
	0x10, 0x21, 0x0C, 0x3A, 0x05, 0x12, 0x56, 0x5B, 0x32, 0x1D, 0x2F, 0x59,
	0x3E, 0x33, 0x2A, 0x2B, 0x26, 0x5E, 0x36, 0x23, 0x17, 0x19, 0x02, 0x28,
	0x1C, 0x2D, 0x04, 0x12, 0x20, 0x00, 0x19, 0x08, 0x05, 0x34, 0x1E, 0x55,
	0x5E, 0x53, 0x6D, 0x2F, 0x59, 0x5D, 0x59, 0x76, 0x09, 0x25, 0x27, 0x5A,
	0x05, 0x1A, 0x56, 0x0B, 0x21, 0x09, 0x5A, 0x59, 0x24, 0x5F, 0x15, 0x09,
	0x15, 0x14, 0x5A, 0x6D, 0x1E, 0x03, 0x07, 0x1A, 0x01, 0x5B, 0x07, 0x45,
	0x12, 0x0C, 0x43, 0x33, 0x1B, 0x13, 0x76, 0x0F, 0x04, 0x57, 0x22, 0x0C,
	0x54, 0x33, 0x29, 0x19, 0x74, 0x1E, 0x38, 0x3B, 0x0F, 0x25, 0x54, 0x07,
	0x39, 0x5F, 0x2C, 0x2B, 0x06, 0x0B, 0x29, 0x2F, 0x2F, 0x26, 0x05, 0x3C,
	0x08, 0x1E, 0x28, 0x3F, 0x09, 0x16, 0x1C, 0x56, 0x2A, 0x40, 0x0E, 0x0B,
	0x39, 0x0C, 0x5A, 0x31, 0x25, 0x27, 0x56, 0x24, 0x28, 0x34, 0x29, 0x27,
	0x05, 0x38, 0x05, 0x37, 0x1F, 0x52, 0x26, 0x05, 0x08, 0x19, 0x25, 0x6D,
	0x00, 0x23, 0x39, 0x2F, 0x24, 0x03, 0x17, 0x07, 0x5F, 0x70, 0x19, 0x19,
	0x0B, 0x02, 0x2C, 0x39, 0x22, 0x02, 0x2A, 0x26, 0x1B, 0x34, 0x0F, 0x5C,
	0x05, 0x04, 0x11, 0x00, 0x01, 0x06, 0x20, 0x13, 0x0A, 0x32, 0x12, 0x28,
	0x53, 0x07, 0x31, 0x15, 0x16, 0x55, 0x20, 0x18, 0x3B, 0x29, 0x02, 0x0D,
	0x24, 0x0D, 0x09, 0x39, 0x2A, 0x12, 0x0A, 0x26, 0x06, 0x00, 0x31, 0x0F,
	0x29, 0x0C, 0x05, 0x1A, 0x27, 0x5F, 0x59, 0x29, 0x44, 0x3A, 0x5B, 0x02,
	0x36, 0x5E, 0x06, 0x0A, 0x54, 0x06, 0x28, 0x24, 0x2F, 0x15, 0x25, 0x1E,
	0x27, 0x35, 0x26, 0x56, 0x33, 0x1A, 0x1F, 0x12, 0x39, 0x3F, 0x7B, 0x1A,
	0x37, 0x2D, 0x29, 0x6D, 0x06, 0x34, 0x59, 0x31, 0x77, 0x0A, 0x52, 0x37,
	0x2A, 0x25, 0x39, 0x2D, 0x1A, 0x07, 0x04, 0x09, 0x06, 0x01, 0x0D, 0x0A,
	0x23, 0x22, 0x1E, 0x5C, 0x09, 0x23, 0x3B, 0x36, 0x22, 0x00, 0x38, 0x12,
	0x5A, 0x07, 0x0C, 0x0E, 0x34, 0x39, 0x5C, 0x08, 0x04, 0x19, 0x5D, 0x12,
	0x0B, 0x3B, 0x50, 0x0F, 0x26, 0x36, 0x07, 0x2D, 0x25, 0x0A, 0x18, 0x1E,
	0x52, 0x01, 0x1B, 0x73, 0x1D, 0x51, 0x18, 0x44, 0x2D, 0x5F, 0x02, 0x1C,
	0x31, 0x6D, 0x14, 0x04, 0x3C, 0x2C, 0x29, 0x1D, 0x14, 0x3C, 0x5A, 0x18,
	0x19, 0x30, 0x3E, 0x33, 0x36, 0x27, 0x00, 0x25, 0x07, 0x74, 0x20, 0x4A,
	0x3E, 0x29, 0x14, 0x2F, 0x26, 0x09, 0x31, 0x28, 0x08, 0x00, 0x5C, 0x5E,
	0x33, 0x34, 0x58, 0x01, 0x13, 0x76, 0x5C, 0x50, 0x3C, 0x11, 0x70, 0x22,
	0x57, 0x36, 0x38, 0x70, 0x1F, 0x17, 0x23, 0x20, 0x23, 0x3F, 0x10, 0x1E,
	0x29, 0x3B, 0x1F, 0x31, 0x3F, 0x05, 0x7B, 0x1A, 0x26, 0x27, 0x27, 0x72,
	0x08, 0x18, 0x0C, 0x3A, 0x37, 0x58, 0x08, 0x0B, 0x13, 0x34, 0x5D, 0x52,
	0x3B, 0x1B, 0x05, 0x2E, 0x51, 0x2C, 0x0A, 0x70, 0x34, 0x05, 0x5B, 0x25,
	0x0B, 0x1F, 0x11, 0x38, 0x5B, 0x2B, 0x3C, 0x11, 0x23, 0x07, 0x2B, 0x36,
	0x34, 0x2D, 0x2E, 0x21, 0x1F, 0x39, 0x0C, 0x02, 0x07, 0x28, 0x59, 0x17,
	0x33, 0x70, 0x59, 0x18, 0x05, 0x23, 0x21, 0x06, 0x2C, 0x45, 0x1B, 0x01,
	0x2D, 0x38, 0x08, 0x12, 0x21, 0x26, 0x35, 0x27, 0x38, 0x33, 0x20, 0x0F,
	0x1E, 0x00, 0x35, 0x3F, 0x10, 0x19, 0x5F, 0x23, 0x08, 0x2C, 0x1F, 0x40,
	0x2C, 0x5A, 0x33, 0x23, 0x2D, 0x33, 0x1F, 0x53, 0x16, 0x12, 0x28, 0x3C,
	0x4E, 0x2D, 0x38, 0x2E, 0x39, 0x00, 0x16, 0x0A, 0x05, 0x5A, 0x31, 0x56,
	0x5F, 0x11, 0x0F, 0x11, 0x3A, 0x3C, 0x17, 0x20, 0x08, 0x0B, 0x19, 0x72,
	0x38, 0x50, 0x25, 0x07, 0x2E, 0x21, 0x51, 0x09, 0x1A, 0x36, 0x5A, 0x07,
	0x1E, 0x2E, 0x2D, 0x18, 0x12, 0x16, 0x29, 0x14, 0x38, 0x18, 0x24, 0x3D,
	0x26, 0x03, 0x39, 0x3F, 0x09, 0x36, 0x5C, 0x3B, 0x01, 0x53, 0x32, 0x1E,
	0x05, 0x17, 0x01, 0x70, 0x27, 0x2C, 0x59, 0x38, 0x20, 0x01, 0x19, 0x5E,
	0x12, 0x36, 0x19, 0x05, 0x5F, 0x00, 0x23, 0x24, 0x20, 0x25, 0x3F, 0x36,
	0x5F, 0x0A, 0x2C, 0x38, 0x31, 0x16, 0x29, 0x1C, 0x28, 0x2D, 0x0A, 0x18,
	0x07, 0x59, 0x10, 0x2D, 0x25, 0x03, 0x1F, 0x13, 0x00, 0x23, 0x57, 0x2E,
	0x70, 0x0D, 0x19, 0x23, 0x38, 0x71, 0x25, 0x0E, 0x04, 0x13, 0x25, 0x20,
	0x0D, 0x29, 0x00, 0x2F, 0x5A, 0x29, 0x0D, 0x1B, 0x72, 0x1E, 0x2E, 0x3F,
	0x09, 0x04, 0x2A, 0x2B, 0x01, 0x20, 0x2A, 0x07, 0x14, 0x41, 0x0A, 0x34,
	0x39, 0x56, 0x26, 0x59, 0x00, 0x55, 0x24, 0x58, 0x3F, 0x21, 0x02, 0x55,
	0x2B, 0x40, 0x29, 0x3C, 0x35, 0x24, 0x12, 0x2B, 0x20, 0x24, 0x3B, 0x03,
	0x15, 0x55, 0x51, 0x21, 0x0C, 0x2E, 0x39, 0x39, 0x1E, 0x1C, 0x1A, 0x27,
	0x17, 0x57, 0x29, 0x14, 0x1A, 0x0D, 0x3E, 0x0E, 0x11, 0x58, 0x28, 0x38,
	0x29, 0x11, 0x5C, 0x0F, 0x36, 0x29, 0x21, 0x5C, 0x0C, 0x57, 0x1A, 0x69,
	0x05, 0x16, 0x0C, 0x3D, 0x20, 0x2D, 0x02, 0x01, 0x1E, 0x23, 0x2F, 0x03,
	0x21, 0x29, 0x10, 0x06, 0x22, 0x1A, 0x1A, 0x23, 0x23, 0x14, 0x38, 0x22,
	0x25, 0x34, 0x18, 0x03, 0x0A, 0x75, 0x0A, 0x35, 0x5C, 0x02, 0x73, 0x06,
	0x12, 0x18, 0x32, 0x04, 0x2D, 0x3B, 0x3D, 0x1F, 0x13, 0x09, 0x50, 0x07,
	0x00, 0x09, 0x08, 0x04, 0x0A, 0x32, 0x30, 0x28, 0x14, 0x06, 0x33, 0x2F,
	0x16, 0x29, 0x07, 0x39, 0x09, 0x5A, 0x51, 0x3F, 0x20, 0x25, 0x18, 0x20,
	0x17, 0x2E, 0x06, 0x34, 0x2E, 0x2F, 0x38, 0x26, 0x35, 0x0C, 0x17, 0x40,
	0x09, 0x02, 0x11, 0x22, 0x3E, 0x16, 0x34, 0x18, 0x3C, 0x04, 0x07, 0x00,
	0x03, 0x01, 0x08, 0x08, 0x22, 0x25, 0x16, 0x0F, 0x08, 0x27, 0x54, 0x0F,
	0x28, 0x38, 0x22, 0x15, 0x06, 0x5C, 0x0B, 0x58, 0x08, 0x09, 0x3B, 0x73,
	0x2E, 0x23, 0x14, 0x28, 0x33, 0x43, 0x25, 0x23, 0x39, 0x03, 0x2A, 0x2E,
	0x23, 0x05, 0x0C, 0x27, 0x29, 0x3B, 0x00, 0x05, 0x08, 0x59, 0x00, 0x2E,
	0x15, 0x47, 0x25, 0x26, 0x5B, 0x20, 0x34, 0x29, 0x59, 0x39, 0x6D, 0x5F,
	0x32, 0x5D, 0x0C, 0x33, 0x2B, 0x2F, 0x5E, 0x2F, 0x1A, 0x3F, 0x03, 0x18,
	0x3B, 0x76, 0x47, 0x0C, 0x09, 0x1D, 0x18, 0x55, 0x28, 0x08, 0x3A, 0x3A,
	0x39, 0x37, 0x03, 0x29, 0x0E, 0x1A, 0x25, 0x28, 0x25, 0x38, 0x5A, 0x02,
	0x25, 0x3C, 0x75, 0x21, 0x18, 0x26, 0x2F, 0x29, 0x0D, 0x1B, 0x04, 0x2C,
	0x06, 0x47, 0x06, 0x41, 0x1E, 0x32, 0x59, 0x07, 0x3B, 0x2A, 0x1A, 0x5A,
	0x53, 0x3D, 0x2F, 0x21, 0x1E, 0x0A, 0x2C, 0x44, 0x72, 0x2D, 0x53, 0x34,
	0x12, 0x0D, 0x34, 0x2D, 0x5D, 0x3B, 0x73, 0x0F, 0x0B, 0x1C, 0x1D, 0x36,
	0x38, 0x2A, 0x57, 0x5A, 0x34, 0x25, 0x2E, 0x56, 0x19, 0x37, 0x34, 0x06,
	0x58, 0x03, 0x3A, 0x1D, 0x0A, 0x0B, 0x19, 0x0C, 0x2F, 0x36, 0x3C, 0x44,
	0x08, 0x06, 0x28, 0x04, 0x00, 0x11, 0x2B, 0x19, 0x0A, 0x03, 0x13, 0x2B,
	0x15, 0x09, 0x0A, 0x17, 0x3D, 0x4A, 0x1E, 0x07, 0x01, 0x3B, 0x33, 0x34,
	0x3C, 0x04, 0x1E, 0x32, 0x34, 0x39, 0x72, 0x5C, 0x28, 0x0A, 0x2D, 0x23,
	0x0B, 0x2A, 0x16, 0x2A, 0x69, 0x39, 0x52, 0x3B, 0x18, 0x27, 0x2D, 0x25,
	0x38, 0x06, 0x71, 0x28, 0x0E, 0x21, 0x5C, 0x26, 0x38, 0x09, 0x06, 0x2D,
	0x30, 0x21, 0x05, 0x3C, 0x23, 0x71, 0x21, 0x56, 0x28, 0x3B, 0x27, 0x3D,
	0x00, 0x17, 0x0C, 0x31, 0x43, 0x4A, 0x59, 0x08, 0x69, 0x09, 0x2A, 0x0F,
	0x06, 0x76, 0x5D, 0x12, 0x1C, 0x33, 0x17, 0x5E, 0x08, 0x3E, 0x05, 0x7B,
	0x22, 0x20, 0x59, 0x0F, 0x74, 0x20, 0x58, 0x58, 0x1F, 0x04, 0x21, 0x4A,
	0x36, 0x02, 0x10, 0x43, 0x23, 0x58, 0x12, 0x73, 0x34, 0x33, 0x57, 0x5B,
	0x17, 0x29, 0x59, 0x58, 0x1C, 0x1A, 0x3F, 0x12, 0x2A, 0x13, 0x32, 0x03,
	0x0F, 0x23, 0x21, 0x35, 0x47, 0x04, 0x5B, 0x08, 0x0D, 0x1B, 0x0E, 0x17,
	0x1F, 0x7B, 0x23, 0x57, 0x5D, 0x1C, 0x70, 0x43, 0x05, 0x1A, 0x0D, 0x0D,
	0x1E, 0x58, 0x05, 0x5F, 0x31, 0x1A, 0x2C, 0x01, 0x5D, 0x04, 0x5D, 0x39,
	0x21, 0x40, 0x11, 0x16, 0x05, 0x08, 0x3B, 0x7B, 0x3B, 0x0A, 0x57, 0x3B,
	0x35, 0x02, 0x54, 0x18, 0x3E, 0x21, 0x07, 0x53, 0x17, 0x20, 0x7A, 0x3E,
	0x26, 0x2F, 0x52, 0x2F, 0x43, 0x32, 0x26, 0x0C, 0x34, 0x3E, 0x35, 0x09,
	0x1D, 0x26, 0x3E, 0x22, 0x34, 0x3E, 0x08, 0x5A, 0x0F, 0x3E, 0x1F, 0x21,
	0x26, 0x3B, 0x57, 0x04, 0x77, 0x19, 0x4A, 0x07, 0x3E, 0x24, 0x3E, 0x56,
	0x07, 0x26, 0x1B, 0x0E, 0x2A, 0x20, 0x13, 0x1A, 0x34, 0x0E, 0x1C, 0x05,
	0x0B, 0x22, 0x56, 0x18, 0x04, 0x31, 0x5F, 0x15, 0x1D, 0x06, 0x13, 0x3D,
	0x17, 0x5B, 0x20, 0x3B, 0x3D, 0x29, 0x09, 0x0D, 0x33, 0x5E, 0x0E, 0x3A,
	0x5A, 0x14, 0x1C, 0x25, 0x25, 0x00, 0x72, 0x06, 0x57, 0x2D, 0x53, 0x08,
	0x2A, 0x37, 0x5E, 0x38, 0x17, 0x3F, 0x53, 0x57, 0x0D, 0x16, 0x25, 0x00,
	0x16, 0x08, 0x23, 0x29, 0x12, 0x39, 0x5F, 0x3B, 0x06, 0x2B, 0x5F, 0x01,
	0x32, 0x05, 0x17, 0x34, 0x18, 0x34, 0x3A, 0x35, 0x1D, 0x0D, 0x2D, 0x03,
	0x04, 0x3A, 0x25, 0x25, 0x5B, 0x32, 0x06, 0x1D, 0x03, 0x1B, 0x51, 0x27,
	0x19, 0x7B, 0x1B, 0x23, 0x21, 0x02, 0x18, 0x5F, 0x0A, 0x3A, 0x22, 0x2F,
	0x08, 0x19, 0x5D, 0x20, 0x30, 0x5A, 0x2D, 0x21, 0x44, 0x07, 0x43, 0x27,
	0x0F, 0x09, 0x0C, 0x25, 0x52, 0x0C, 0x25, 0x32, 0x3A, 0x4E, 0x3D, 0x1C,
	0x36, 0x3E, 0x17, 0x1F, 0x2C, 0x03, 0x21, 0x26, 0x00, 0x21, 0x0F, 0x02,
	0x0E, 0x1A, 0x23, 0x09, 0x5C, 0x53, 0x14, 0x2A, 0x74, 0x35, 0x37, 0x0D,
	0x25, 0x69, 0x2F, 0x10, 0x05, 0x23, 0x32, 0x5F, 0x28, 0x0B, 0x32, 0x2F,
	0x1E, 0x39, 0x57, 0x0C, 0x33, 0x0A, 0x54, 0x26, 0x2F, 0x70, 0x5B, 0x13,
	0x1A, 0x40, 0x34, 0x0A, 0x05, 0x45, 0x39, 0x71, 0x05, 0x0C, 0x1A, 0x24,
	0x76, 0x58, 0x34, 0x34, 0x38, 0x31, 0x36, 0x0D, 0x3A, 0x1A, 0x17, 0x2D,
	0x4A, 0x5B, 0x27, 0x29, 0x02, 0x4E, 0x1C, 0x1B, 0x26, 0x39, 0x0A, 0x29,
	0x5D, 0x3B, 0x24, 0x0E, 0x1A, 0x06, 0x77, 0x00, 0x22, 0x07, 0x05, 0x3A,
	0x09, 0x04, 0x5D, 0x3F, 0x6D, 0x21, 0x56, 0x1C, 0x0D, 0x73, 0x2F, 0x2C,
	0x28, 0x08, 0x0E, 0x19, 0x00, 0x38, 0x5A, 0x1A, 0x34, 0x18, 0x56, 0x58,
	0x23, 0x08, 0x17, 0x3F, 0x5F, 0x2D, 0x26, 0x24, 0x1F, 0x23, 0x18, 0x1E,
	0x25, 0x14, 0x5F, 0x11, 0x02, 0x58, 0x5C, 0x2A, 0x28, 0x5A, 0x23, 0x45,
	0x02, 0x14, 0x39, 0x18, 0x0A, 0x2C, 0x18, 0x08, 0x23, 0x3B, 0x25, 0x75,
	0x34, 0x4A, 0x5F, 0x03, 0x35, 0x2D, 0x53, 0x5E, 0x19, 0x24, 0x5E, 0x19,
	0x1F, 0x11, 0x7A, 0x5B, 0x29, 0x5F, 0x2F, 0x0C, 0x1F, 0x03, 0x05, 0x33,
	0x1A, 0x3D, 0x18, 0x58, 0x00, 0x08, 0x20, 0x27, 0x17, 0x1F, 0x15, 0x05,
	0x53, 0x22, 0x3E, 0x1B, 0x34, 0x57, 0x22, 0x44, 0x05, 0x2B, 0x30, 0x2C,
	0x24, 0x7B, 0x38, 0x0D, 0x3F, 0x04, 0x26, 0x5F, 0x08, 0x57, 0x2F, 0x12,
	0x09, 0x05, 0x37, 0x3B, 0x2C, 0x0F, 0x13, 0x57, 0x5A, 0x69, 0x1C, 0x59,
	0x3C, 0x1D, 0x21, 0x1F, 0x20, 0x0D, 0x5A, 0x31, 0x01, 0x06, 0x02, 0x22,
	0x25, 0x03, 0x00, 0x09, 0x59, 0x0D, 0x5F, 0x31, 0x1A, 0x3F, 0x30, 0x00,
	0x4E, 0x39, 0x5C, 0x77, 0x2B, 0x4A, 0x04, 0x2F, 0x0A, 0x5A, 0x27, 0x03,
	0x2A, 0x30, 0x55, 0x29, 0x01, 0x08, 0x33, 0x43, 0x30, 0x5F, 0x5F, 0x06,
	0x0A, 0x38, 0x38, 0x5F, 0x38, 0x3B, 0x0F, 0x38, 0x0F, 0x09, 0x3B, 0x27,
	0x38, 0x21, 0x15, 0x06, 0x09, 0x37, 0x1B, 0x75, 0x07, 0x0A, 0x26, 0x40,
	0x0F, 0x22, 0x03, 0x1A, 0x05, 0x16, 0x04, 0x06, 0x28, 0x18, 0x03, 0x54,
	0x1B, 0x0A, 0x1A, 0x2F, 0x2F, 0x35, 0x57, 0x0C, 0x38, 0x1D, 0x08, 0x3C,
	0x5E, 0x70, 0x28, 0x2E, 0x5B, 0x25, 0x70, 0x0B, 0x38, 0x39, 0x1E, 0x05,
	0x5B, 0x1B, 0x29, 0x3E, 0x11, 0x03, 0x24, 0x0C, 0x06, 0x2D, 0x58, 0x26,
	0x2D, 0x11, 0x75, 0x47, 0x25, 0x14, 0x04, 0x32, 0x23, 0x0A, 0x22, 0x0E,
	0x6D, 0x1D, 0x24, 0x36, 0x0A, 0x70, 0x55, 0x53, 0x01, 0x5C, 0x69, 0x0D,
	0x09, 0x07, 0x11, 0x7A, 0x03, 0x27, 0x17, 0x3D, 0x2B, 0x5E, 0x03, 0x24,
	0x5D, 0x2C, 0x18, 0x32, 0x1C, 0x2E, 0x0E, 0x27, 0x2D, 0x5D, 0x2F, 0x74,
	0x3B, 0x00, 0x2C, 0x2F, 0x73, 0x1D, 0x22, 0x34, 0x23, 0x0D, 0x55, 0x06,
	0x04, 0x3C, 0x2F, 0x58, 0x05, 0x1F, 0x5F, 0x6D, 0x24, 0x14, 0x01, 0x02,
	0x34, 0x5E, 0x56, 0x25, 0x5E, 0x2E, 0x16, 0x51, 0x2D, 0x0F, 0x0C, 0x1B,
	0x20, 0x08, 0x1C, 0x77, 0x47, 0x33, 0x01, 0x26, 0x32, 0x5C, 0x0C, 0x18,
	0x28, 0x76, 0x0D, 0x36, 0x1F, 0x07, 0x35, 0x54, 0x18, 0x34, 0x3F, 0x23,
	0x04, 0x59, 0x02, 0x3D, 0x77, 0x3B, 0x28, 0x22, 0x1C, 0x6D, 0x2F, 0x57,
	0x45, 0x58, 0x15, 0x2E, 0x28, 0x2C, 0x5F, 0x35, 0x1B, 0x00, 0x5E, 0x3B,
	0x27, 0x2B, 0x35, 0x29, 0x1A, 0x23, 0x0D, 0x35, 0x29, 0x12, 0x2A, 0x23,
	0x07, 0x3B, 0x20, 0x21, 0x3A, 0x50, 0x03, 0x08, 0x06, 0x34, 0x10, 0x0D,
	0x24, 0x2A, 0x36, 0x0F, 0x3E, 0x01, 0x35, 0x2B, 0x36, 0x24, 0x1C, 0x26,
	0x2B, 0x52, 0x2C, 0x0F, 0x3A, 0x59, 0x50, 0x0C, 0x02, 0x33, 0x55, 0x25,
	0x04, 0x23, 0x2D, 0x00, 0x34, 0x07, 0x1D, 0x30, 0x5E, 0x20, 0x0D, 0x03,
	0x05, 0x2E, 0x50, 0x45, 0x1A, 0x33, 0x59, 0x0A, 0x2F, 0x31, 0x15, 0x1A,
	0x3B, 0x0A, 0x0C, 0x11, 0x1C, 0x36, 0x1C, 0x05, 0x36, 0x09, 0x09, 0x23,
	0x5F, 0x37, 0x14, 0x12, 0x5D, 0x5C, 0x06, 0x04, 0x19, 0x59, 0x22, 0x7B,
	0x47, 0x0F, 0x3B, 0x53, 0x7A, 0x1E, 0x22, 0x21, 0x5E, 0x14, 0x34, 0x31,
	0x18, 0x01, 0x1B, 0x38, 0x07, 0x34, 0x3C, 0x00, 0x38, 0x2F, 0x3A, 0x2C,
	0x7B, 0x26, 0x57, 0x59, 0x2C, 0x29, 0x5A, 0x4E, 0x57, 0x06, 0x12, 0x1C,
	0x15, 0x39, 0x58, 0x03, 0x55, 0x2F, 0x37, 0x3B, 0x16, 0x27, 0x59, 0x22,
	0x3C, 0x72, 0x3B, 0x3B, 0x26, 0x1B, 0x70, 0x1C, 0x3B, 0x2F, 0x11, 0x16,
	0x19, 0x10, 0x2C, 0x1A, 0x73, 0x35, 0x56, 0x00, 0x2F, 0x0D, 0x0A, 0x2C,
	0x58, 0x2E, 0x31, 0x43, 0x0C, 0x18, 0x2A, 0x3B, 0x3F, 0x0F, 0x04, 0x5A,
	0x25, 0x25, 0x30, 0x06, 0x1C, 0x36, 0x23, 0x17, 0x2D, 0x32, 0x29, 0x5D,
	0x2E, 0x1B, 0x0D, 0x31, 0x19, 0x10, 0x5A, 0x01, 0x0A, 0x00, 0x09, 0x26,
	0x25, 0x23, 0x1A, 0x58, 0x34, 0x0A, 0x06, 0x43, 0x1B, 0x5A, 0x23, 0x30,
	0x22, 0x03, 0x1D, 0x1B, 0x74, 0x3E, 0x23, 0x0A, 0x23, 0x34, 0x35, 0x11,
	0x45, 0x1D, 0x24, 0x2A, 0x52, 0x3F, 0x18, 0x72, 0x1F, 0x26, 0x28, 0x33,
	0x24, 0x15, 0x15, 0x36, 0x18, 0x77, 0x00, 0x53, 0x08, 0x3F, 0x2C, 0x47,
	0x07, 0x3C, 0x0E, 0x34, 0x2E, 0x59, 0x56, 0x27, 0x20, 0x2F, 0x11, 0x2F,
	0x27, 0x2F, 0x03, 0x55, 0x06, 0x02, 0x0E, 0x47, 0x07, 0x3A, 0x31, 0x00,
	0x16, 0x27, 0x02, 0x1C, 0x06, 0x0E, 0x0E, 0x2D, 0x1E, 0x27, 0x07, 0x00,
	0x57, 0x22, 0x35, 0x59, 0x18, 0x00, 0x26, 0x0C, 0x38, 0x09, 0x08, 0x0A,
	0x3A, 0x38, 0x39, 0x04, 0x3E, 0x7B, 0x02, 0x0A, 0x5C, 0x04, 0x09, 0x1E,
	0x2A, 0x2D, 0x3E, 0x35, 0x08, 0x13, 0x0A, 0x21, 0x11, 0x04, 0x0F, 0x0B,
	0x27, 0x1A, 0x5E, 0x02, 0x3C, 0x05, 0x71, 0x59, 0x23, 0x25, 0x5D, 0x7B,
	0x38, 0x29, 0x2A, 0x02, 0x37, 0x24, 0x0F, 0x3D, 0x22, 0x11, 0x58, 0x53,
	0x24, 0x04, 0x36, 0x3B, 0x38, 0x2D, 0x3B, 0x14, 0x22, 0x19, 0x5D, 0x5C,
	0x08, 0x2D, 0x32, 0x58, 0x07, 0x00, 0x19, 0x35, 0x17, 0x2C, 0x2E, 0x5F,
	0x24, 0x5D, 0x1E, 0x3A, 0x23, 0x2E, 0x28, 0x2D, 0x04, 0x2A, 0x56, 0x09,
	0x58, 0x27, 0x55, 0x18, 0x2D, 0x58, 0x34, 0x5F, 0x32, 0x5D, 0x04, 0x0A,
	0x15, 0x03, 0x02, 0x2A, 0x30, 0x43, 0x25, 0x5C, 0x28, 0x0D, 0x20, 0x2A,
	0x26, 0x07, 0x0E, 0x34, 0x04, 0x58, 0x5F, 0x16, 0x3A, 0x4E, 0x5C, 0x08,
	0x32, 0x01, 0x57, 0x0F, 0x3A, 0x0A, 0x0A, 0x20, 0x17, 0x28, 0x2E, 0x5C,
	0x22, 0x09, 0x2E, 0x3B, 0x1A, 0x32, 0x5A, 0x0D, 0x32, 0x07, 0x2D, 0x5F,
	0x5D, 0x24, 0x5B, 0x15, 0x0C, 0x11, 0x71, 0x1B, 0x11, 0x58, 0x5E, 0x29,
	0x01, 0x23, 0x1D, 0x52, 0x2A, 0x2D, 0x27, 0x0A, 0x0E, 0x7B, 0x5E, 0x0B,
	0x3A, 0x5B, 0x06, 0x47, 0x30, 0x04, 0x2F, 0x3A, 0x19, 0x33, 0x23, 0x2F,
	0x25, 0x03, 0x04, 0x1B, 0x2A, 0x15, 0x3A, 0x35, 0x38, 0x28, 0x18, 0x05,
	0x2A, 0x3D, 0x2F, 0x24, 0x58, 0x0A, 0x0F, 0x01, 0x76, 0x21, 0x19, 0x18,
	0x07, 0x27, 0x3F, 0x27, 0x1B, 0x3F, 0x1B, 0x35, 0x30, 0x1E, 0x18, 0x0E,
	0x54, 0x0A, 0x59, 0x21, 0x07, 0x3B, 0x51, 0x45, 0x18, 0x72, 0x47, 0x22,
	0x17, 0x05, 0x16, 0x2F, 0x23, 0x2B, 0x05, 0x21, 0x1C, 0x27, 0x5A, 0x25,
	0x05, 0x0B, 0x37, 0x39, 0x1B, 0x35, 0x5D, 0x10, 0x1D, 0x39, 0x32, 0x1E,
	0x24, 0x08, 0x3A, 0x09, 0x18, 0x20, 0x1D, 0x33, 0x2C, 0x1B, 0x03, 0x28,
	0x58, 0x2B, 0x00, 0x14, 0x59, 0x20, 0x75, 0x39, 0x2B, 0x1B, 0x2D, 0x2A,
	0x34, 0x33, 0x41, 0x0A, 0x30, 0x28, 0x0E, 0x36, 0x09, 0x0F, 0x3C, 0x54,
	0x39, 0x3D, 0x76, 0x2D, 0x12, 0x04, 0x3E, 0x73, 0x24, 0x57, 0x0A, 0x07,
	0x70, 0x00, 0x23, 0x18, 0x3F, 0x75, 0x20, 0x55, 0x37, 0x0C, 0x06, 0x5C,
	0x26, 0x56, 0x0E, 0x01, 0x25, 0x2B, 0x1B, 0x0D, 0x20, 0x3F, 0x4A, 0x3F,
	0x3B, 0x75, 0x3E, 0x14, 0x06, 0x5F, 0x35, 0x23, 0x20, 0x3C, 0x20, 0x23,
	0x02, 0x1B, 0x00, 0x25, 0x28, 0x5C, 0x06, 0x02, 0x24, 0x14, 0x5E, 0x35,
	0x05, 0x5C, 0x01, 0x07, 0x34, 0x0F, 0x09, 0x0E, 0x5C, 0x52, 0x09, 0x1D,
	0x32, 0x3F, 0x20, 0x22, 0x1F, 0x07, 0x1E, 0x2A, 0x3F, 0x03, 0x28, 0x05,
	0x12, 0x24, 0x31, 0x26, 0x15, 0x0E, 0x20, 0x26, 0x36, 0x59, 0x30, 0x3E,
	0x3E, 0x1B, 0x3B, 0x56, 0x1C, 0x33, 0x72, 0x02, 0x0E, 0x0D, 0x1B, 0x2A,
	0x05, 0x25, 0x04, 0x24, 0x09, 0x02, 0x25, 0x01, 0x1F, 0x03, 0x2B, 0x50,
	0x08, 0x04, 0x28, 0x3B, 0x26, 0x45, 0x21, 0x14, 0x43, 0x54, 0x5F, 0x2F,
	0x24, 0x5C, 0x15, 0x18, 0x01, 0x31, 0x09, 0x13, 0x41, 0x33, 0x12, 0x24,
	0x06, 0x29, 0x19, 0x12, 0x29, 0x37, 0x0A, 0x1F, 0x10, 0x59, 0x3B, 0x1F,
	0x02, 0x0A, 0x07, 0x59, 0x0A, 0x08, 0x31, 0x3E, 0x50, 0x58, 0x0A, 0x24,
	0x5A, 0x07, 0x57, 0x1C, 0x30, 0x19, 0x0B, 0x25, 0x09, 0x3A, 0x3F, 0x58,
	0x25, 0x09, 0x10, 0x16, 0x59, 0x39, 0x02, 0x37, 0x14, 0x37, 0x2C, 0x40,
	0x33, 0x1B, 0x30, 0x0F, 0x3E, 0x7B, 0x58, 0x11, 0x1F, 0x3C, 0x31, 0x43,
	0x02, 0x25, 0x2F, 0x29, 0x5B, 0x07, 0x09, 0x29, 0x10, 0x2B, 0x2A, 0x3D,
	0x21, 0x00, 0x15, 0x32, 0x56, 0x05, 0x27, 0x3A, 0x16, 0x56, 0x1C, 0x71,
	0x1C, 0x11, 0x08, 0x3A, 0x71, 0x01, 0x38, 0x27, 0x2F, 0x72, 0x3F, 0x09,
	0x06, 0x58, 0x35, 0x5E, 0x08, 0x3B, 0x04, 0x33, 0x15, 0x15, 0x45, 0x5C,
	0x7B, 0x2B, 0x23, 0x2C, 0x44, 0x29, 0x0F, 0x16, 0x06, 0x3C, 0x28, 0x23,
	0x2E, 0x19, 0x3C, 0x33, 0x00, 0x58, 0x37, 0x03, 0x3A, 0x3C, 0x1B, 0x5B,
	0x5F, 0x05, 0x29, 0x34, 0x3E, 0x0F, 0x29, 0x3D, 0x32, 0x5F, 0x0A, 0x04,
	0x36, 0x23, 0x1B, 0x07, 0x6D, 0x2A, 0x0C, 0x5B, 0x00, 0x7A, 0x1A, 0x29,
	0x3D, 0x23, 0x09, 0x06, 0x07, 0x1A, 0x5D, 0x15, 0x5C, 0x0B, 0x5E, 0x5C,
	0x70, 0x3B, 0x4A, 0x0A, 0x40, 0x10, 0x55, 0x2B, 0x5D, 0x18, 0x69, 0x05,
	0x13, 0x00, 0x0D, 0x2B, 0x5F, 0x17, 0x00, 0x07, 0x1A, 0x1E, 0x1B, 0x02,
	0x28, 0x28, 0x09, 0x53, 0x01, 0x08, 0x0C, 0x5C, 0x29, 0x37, 0x28, 0x32,
	0x20, 0x05, 0x18, 0x26, 0x16, 0x15, 0x2B, 0x26, 0x44, 0x11, 0x1B, 0x2C,
	0x2B, 0x26, 0x3B, 0x2D, 0x18, 0x3F, 0x09, 0x2B, 0x27, 0x0B, 0x37, 0x0D,
	0x35, 0x3B, 0x15, 0x0D, 0x3B, 0x70, 0x35, 0x34, 0x36, 0x5A, 0x0E, 0x05,
	0x14, 0x2D, 0x40, 0x29, 0x26, 0x38, 0x29, 0x3C, 0x07, 0x29, 0x59, 0x26,
	0x3C, 0x05, 0x07, 0x0F, 0x3E, 0x25, 0x01, 0x26, 0x08, 0x5E, 0x5F, 0x0B,
	0x0E, 0x00, 0x21, 0x3E, 0x0C, 0x29, 0x16, 0x24, 0x38, 0x14, 0x5F, 0x54,
	0x5C, 0x5E, 0x20, 0x39, 0x51, 0x59, 0x3E, 0x27, 0x54, 0x34, 0x57, 0x01,
	0x27, 0x35, 0x32, 0x57, 0x00, 0x2F, 0x26, 0x02, 0x3D, 0x5C, 0x27, 0x0F,
	0x36, 0x24, 0x18, 0x2E, 0x0E, 0x50, 0x45, 0x0E, 0x1A, 0x34, 0x18, 0x03,
	0x59, 0x24, 0x3A, 0x2E, 0x18, 0x5D, 0x34, 0x36, 0x03, 0x05, 0x04, 0x38,
	0x25, 0x2C, 0x03, 0x0D, 0x17, 0x34, 0x13, 0x26, 0x00, 0x2E, 0x00, 0x57,
	0x17, 0x0A, 0x75, 0x54, 0x0F, 0x1F, 0x3C, 0x6D, 0x5B, 0x2D, 0x0A, 0x33,
	0x35, 0x14, 0x37, 0x02, 0x12, 0x00, 0x3E, 0x2F, 0x38, 0x3F, 0x07, 0x5F,
	0x52, 0x37, 0x06, 0x77, 0x3F, 0x35, 0x5B, 0x33, 0x75, 0x2F, 0x39, 0x0C,
	0x21, 0x11, 0x34, 0x56, 0x04, 0x5E, 0x2A, 0x1A, 0x0E, 0x3C, 0x5A, 0x71,
	0x3D, 0x53, 0x2F, 0x24, 0x13, 0x08, 0x4E, 0x21, 0x58, 0x35, 0x5D, 0x35,
	0x5F, 0x1C, 0x0E, 0x04, 0x51, 0x41, 0x3A, 0x0B, 0x34, 0x10, 0x1D, 0x03,
	0x0C, 0x20, 0x0F, 0x02, 0x18, 0x07, 0x1F, 0x04, 0x03, 0x3D, 0x31, 0x2D,
	0x29, 0x3D, 0x3D, 0x0C, 0x1D, 0x15, 0x17, 0x28, 0x31, 0x03, 0x3B, 0x0C,
	0x25, 0x30, 0x38, 0x0B, 0x03, 0x38, 0x0E, 0x3B, 0x32, 0x02, 0x2A, 0x76,
	0x23, 0x10, 0x08, 0x5E, 0x07, 0x47, 0x51, 0x3C, 0x5C, 0x70, 0x1B, 0x06,
	0x3B, 0x5D, 0x32, 0x27, 0x02, 0x21, 0x38, 0x11, 0x38, 0x1B, 0x07, 0x53,
	0x0A, 0x35, 0x2A, 0x1C, 0x32, 0x17, 0x2F, 0x09, 0x57, 0x5A, 0x0D, 0x04,
	0x0E, 0x3C, 0x27, 0x3A, 0x0F, 0x15, 0x3E, 0x40, 0x20, 0x2B, 0x59, 0x3A,
	0x1D, 0x1B, 0x47, 0x0B, 0x3F, 0x13, 0x1A, 0x25, 0x0B, 0x3F, 0x3C, 0x26,
	0x5D, 0x07, 0x34, 0x33, 0x2E, 0x09, 0x17, 0x57, 0x5E, 0x7B, 0x05, 0x4E,
	0x2D, 0x11, 0x33, 0x3E, 0x29, 0x25, 0x04, 0x07, 0x3E, 0x17, 0x2F, 0x06,
	0x2E, 0x43, 0x16, 0x28, 0x07, 0x0C, 0x16, 0x37, 0x06, 0x1A, 0x70, 0x28,
	0x2F, 0x38, 0x2C, 0x17, 0x5F, 0x16, 0x22, 0x3D, 0x08, 0x28, 0x55, 0x38,
	0x08, 0x0B, 0x14, 0x14, 0x1A, 0x07, 0x21, 0x08, 0x06, 0x0D, 0x19, 0x6D,
	0x03, 0x19, 0x20, 0x06, 0x36, 0x47, 0x2A, 0x58, 0x39, 0x29, 0x07, 0x28,
	0x0B, 0x2D, 0x31, 0x29, 0x57, 0x5F, 0x0A, 0x2D, 0x29, 0x02, 0x08, 0x04,
	0x07, 0x5A, 0x1B, 0x1B, 0x05, 0x12, 0x27, 0x14, 0x0B, 0x2E, 0x0F, 0x01,
	0x2C, 0x45, 0x0E, 0x75, 0x5E, 0x54, 0x0B, 0x53, 0x77, 0x2D, 0x32, 0x02,
	0x1C, 0x1B, 0x26, 0x57, 0x37, 0x03, 0x14, 0x09, 0x39, 0x2D, 0x18, 0x0F,
	0x5B, 0x22, 0x04, 0x09, 0x72, 0x0E, 0x10, 0x06, 0x3B, 0x32, 0x35, 0x37,
	0x2D, 0x39, 0x21, 0x3A, 0x53, 0x1C, 0x0A, 0x75, 0x54, 0x26, 0x25, 0x09,
	0x0E, 0x07, 0x2F, 0x0D, 0x19, 0x76, 0x3C, 0x2C, 0x1B, 0x0E, 0x11, 0x55,
	0x33, 0x08, 0x22, 0x27, 0x58, 0x0C, 0x14, 0x20, 0x05, 0x2F, 0x54, 0x38,
	0x19, 0x21, 0x21, 0x02, 0x04, 0x2C, 0x75, 0x2B, 0x35, 0x2B, 0x2D, 0x37,
	0x34, 0x2F, 0x34, 0x2C, 0x34, 0x29, 0x2C, 0x39, 0x0A, 0x35, 0x25, 0x18,
	0x56, 0x02, 0x29, 0x18, 0x51, 0x39, 0x2A, 0x15, 0x5E, 0x0D, 0x1E, 0x13,
	0x01, 0x16, 0x12, 0x41, 0x18, 0x0E, 0x38, 0x23, 0x3B, 0x0F, 0x04, 0x1E,
	0x16, 0x1F, 0x1C, 0x75, 0x04, 0x25, 0x21, 0x3A, 0x18, 0x3A, 0x35, 0x58,
	0x1A, 0x71, 0x2D, 0x55, 0x19, 0x08, 0x15, 0x19, 0x34, 0x0B, 0x5C, 0x7A,
	0x24, 0x36, 0x25, 0x5A, 0x0A, 0x0D, 0x17, 0x36, 0x0E, 0x73, 0x2D, 0x0E,
	0x29, 0x1C, 0x09, 0x1D, 0x0D, 0x09, 0x5A, 0x17, 0x1E, 0x32, 0x18, 0x5A,
	0x69, 0x5A, 0x15, 0x16, 0x1C, 0x15, 0x18, 0x12, 0x41, 0x44, 0x76, 0x3C,
	0x22, 0x2D, 0x5D, 0x21, 0x2F, 0x2E, 0x28, 0x5D, 0x09, 0x58, 0x09, 0x2A,
	0x2E, 0x04, 0x1A, 0x3B, 0x25, 0x22, 0x24, 0x47, 0x06, 0x29, 0x20, 0x30,
	0x24, 0x12, 0x39, 0x09, 0x72, 0x14, 0x10, 0x37, 0x2A, 0x21, 0x1C, 0x16,
	0x2F, 0x3C, 0x16, 0x29, 0x53, 0x01, 0x1A, 0x1A, 0x1E, 0x0D, 0x17, 0x53,
	0x1B, 0x20, 0x14, 0x1B, 0x33, 0x71, 0x01, 0x50, 0x34, 0x3A, 0x77, 0x1E,
	0x10, 0x41, 0x31, 0x27, 0x38, 0x4A, 0x22, 0x5F, 0x2E, 0x24, 0x05, 0x25,
	0x06, 0x71, 0x1B, 0x0C, 0x3F, 0x09, 0x69, 0x5E, 0x37, 0x5B, 0x1C, 0x3A,
	0x3D, 0x04, 0x05, 0x04, 0x2C, 0x58, 0x51, 0x5E, 0x24, 0x18, 0x00, 0x2F,
	0x08, 0x0C, 0x73, 0x5F, 0x08, 0x28, 0x3C, 0x6D, 0x36, 0x57, 0x57, 0x29,
	0x2F, 0x34, 0x57, 0x25, 0x1E, 0x24, 0x0F, 0x39, 0x58, 0x2A, 0x30, 0x2A,
	0x0C, 0x22, 0x52, 0x2D, 0x07, 0x08, 0x5A, 0x3C, 0x29, 0x18, 0x28, 0x28,
	0x08, 0x2A, 0x55, 0x03, 0x5D, 0x3C, 0x06, 0x47, 0x36, 0x3A, 0x53, 0x76,
	0x07, 0x52, 0x2C, 0x40, 0x14, 0x0E, 0x0A, 0x1E, 0x38, 0x28, 0x38, 0x51,
	0x2D, 0x19, 0x28, 0x20, 0x15, 0x3D, 0x05, 0x0D, 0x2A, 0x0D, 0x5E, 0x0F,
	0x26, 0x2B, 0x39, 0x58, 0x22, 0x27, 0x25, 0x09, 0x2C, 0x2C, 0x70, 0x3F,
	0x1B, 0x05, 0x00, 0x30, 0x22, 0x14, 0x24, 0x59, 0x12, 0x5A, 0x55, 0x25,
	0x2F, 0x31, 0x0A, 0x05, 0x41, 0x2C, 0x6D, 0x5B, 0x57, 0x19, 0x3B, 0x30,
	0x38, 0x2A, 0x16, 0x28, 0x7B, 0x59, 0x2F, 0x58, 0x1D, 0x21, 0x5F, 0x23,
	0x3A, 0x31, 0x1A, 0x01, 0x14, 0x2A, 0x53, 0x00, 0x0D, 0x2B, 0x29, 0x53,
	0x0B, 0x5C, 0x37, 0x17, 0x26, 0x01, 0x47, 0x10, 0x0A, 0x3E, 0x0A, 0x39,
	0x04, 0x1A, 0x3A, 0x12, 0x18, 0x39, 0x41, 0x59, 0x0F, 0x26, 0x52, 0x04,
	0x5B, 0x26, 0x15, 0x56, 0x45, 0x44, 0x15, 0x2F, 0x2B, 0x5F, 0x5F, 0x15,
	0x0F, 0x29, 0x39, 0x53, 0x2F, 0x2D, 0x52, 0x1F, 0x04, 0x0D, 0x43, 0x22,
	0x39, 0x2F, 0x7B, 0x1A, 0x17, 0x39, 0x2A, 0x03, 0x08, 0x39, 0x5E, 0x40,
	0x0E, 0x0F, 0x20, 0x2C, 0x01, 0x24, 0x55, 0x0D, 0x1E, 0x01, 0x12, 0x36,
	0x36, 0x5B, 0x03, 0x70, 0x29, 0x2A, 0x23, 0x2D, 0x71, 0x0F, 0x06, 0x5E,
	0x01, 0x17, 0x5A, 0x31, 0x09, 0x2E, 0x33, 0x28, 0x0C, 0x05, 0x28, 0x0C,
	0x25, 0x34, 0x29, 0x11, 0x17, 0x29, 0x18, 0x41, 0x0D, 0x32, 0x01, 0x11,
	0x2B, 0x27, 0x14, 0x21, 0x09, 0x0C, 0x03, 0x76, 0x0A, 0x03, 0x57, 0x2C,
	0x2D, 0x3E, 0x56, 0x1F, 0x04, 0x20, 0x39, 0x15, 0x07, 0x38, 0x18, 0x38,
	0x57, 0x1B, 0x1A, 0x30, 0x01, 0x29, 0x01, 0x5A, 0x0B, 0x2B, 0x17, 0x26,
	0x33, 0x28, 0x03, 0x56, 0x0F, 0x11, 0x36, 0x09, 0x33, 0x03, 0x33, 0x04,
	0x1E, 0x04, 0x0B, 0x25, 0x1A, 0x21, 0x2A, 0x08, 0x2D, 0x27, 0x43, 0x15,
	0x02, 0x59, 0x0E, 0x36, 0x31, 0x56, 0x5D, 0x2B, 0x35, 0x07, 0x37, 0x0C,
	0x75, 0x1C, 0x2F, 0x0D, 0x3E, 0x20, 0x2A, 0x0E, 0x0A, 0x38, 0x7A, 0x26,
	0x59, 0x0F, 0x22, 0x7A, 0x55, 0x25, 0x25, 0x1B, 0x0D, 0x3C, 0x51, 0x02,
	0x01, 0x00, 0x0A, 0x0A, 0x58, 0x31, 0x21, 0x2B, 0x27, 0x21, 0x3F, 0x15,
	0x00, 0x54, 0x02, 0x1A, 0x04, 0x15, 0x12, 0x1B, 0x2D, 0x27, 0x05, 0x22,
	0x2F, 0x3A, 0x14, 0x5A, 0x2B, 0x5E, 0x53, 0x35, 0x5D, 0x31, 0x3A, 0x11,
	0x05, 0x55, 0x17, 0x1B, 0x18, 0x75, 0x1F, 0x53, 0x16, 0x0D, 0x3A, 0x06,
	0x1B, 0x34, 0x3B, 0x07, 0x59, 0x05, 0x2C, 0x1B, 0x2F, 0x19, 0x0D, 0x0F,
	0x07, 0x00, 0x0E, 0x39, 0x0F, 0x2D, 0x3B, 0x16, 0x14, 0x34, 0x19, 0x18,
	0x0D, 0x06, 0x39, 0x3B, 0x1A, 0x35, 0x4E, 0x26, 0x58, 0x33, 0x0E, 0x32,
	0x1C, 0x06, 0x34, 0x3A, 0x31, 0x19, 0x11, 0x1B, 0x01, 0x08, 0x28, 0x58,
	0x27, 0x1D, 0x23, 0x1D, 0x02, 0x17, 0x19, 0x11, 0x2B, 0x26, 0x28, 0x03,
	0x11, 0x08, 0x1D, 0x33, 0x04, 0x59, 0x37, 0x3D, 0x3B, 0x3B, 0x51, 0x20,
	0x0A, 0x0A, 0x0E, 0x0C, 0x2B, 0x01, 0x26, 0x1C, 0x37, 0x5E, 0x1D, 0x15,
	0x25, 0x2F, 0x5B, 0x1A, 0x31, 0x3C, 0x2C, 0x3F, 0x2F, 0x29, 0x21, 0x56,
	0x19, 0x58, 0x11, 0x14, 0x30, 0x07, 0x58, 0x04, 0x0E, 0x2C, 0x0B, 0x2C,
	0x31, 0x5A, 0x0F, 0x5D, 0x5B, 0x23, 0x3A, 0x20, 0x23, 0x2A, 0x1A, 0x28,
	0x51, 0x36, 0x3D, 0x3B, 0x0A, 0x20, 0x01, 0x06, 0x7B, 0x47, 0x22, 0x21,
	0x09, 0x2E, 0x01, 0x14, 0x3C, 0x39, 0x73, 0x04, 0x24, 0x3B, 0x03, 0x09,
	0x09, 0x56, 0x08, 0x32, 0x13, 0x34, 0x13, 0x29, 0x52, 0x37, 0x55, 0x0E,
	0x04, 0x1D, 0x0F, 0x2B, 0x10, 0x5A, 0x39, 0x20, 0x43, 0x09, 0x24, 0x09,
	0x7A, 0x29, 0x11, 0x5B, 0x02, 0x11, 0x5D, 0x55, 0x00, 0x3E, 0x73, 0x3C,
	0x25, 0x01, 0x5A, 0x24, 0x36, 0x31, 0x3A, 0x06, 0x0D, 0x24, 0x52, 0x08,
	0x33, 0x71, 0x5A, 0x2C, 0x3E, 0x07, 0x05, 0x01, 0x09, 0x02, 0x12, 0x20,
	0x35, 0x0D, 0x27, 0x21, 0x2E, 0x16, 0x23, 0x3C, 0x01, 0x0F, 0x2D, 0x06,
	0x18, 0x0C, 0x0E, 0x5B, 0x39, 0x19, 0x3B, 0x20, 0x5D, 0x13, 0x25, 0x01,
	0x71, 0x19, 0x2E, 0x3F, 0x3C, 0x7B, 0x24, 0x02, 0x07, 0x06, 0x10, 0x59,
	0x2C, 0x1D, 0x0A, 0x09, 0x5C, 0x18, 0x59, 0x0F, 0x30, 0x58, 0x53, 0x20,
	0x13, 0x37, 0x59, 0x31, 0x20, 0x5C, 0x73, 0x35, 0x26, 0x41, 0x1D, 0x7A,
	0x07, 0x4E, 0x1C, 0x05, 0x36, 0x36, 0x29, 0x3C, 0x03, 0x12, 0x34, 0x19,
	0x1D, 0x0C, 0x37, 0x2E, 0x10, 0x2A, 0x39, 0x0D, 0x55, 0x2B, 0x1D, 0x32,
	0x17, 0x3E, 0x04, 0x0A, 0x58, 0x73, 0x22, 0x2C, 0x0D, 0x40, 0x09, 0x1A,
	0x3B, 0x1D, 0x31, 0x27, 0x0A, 0x33, 0x59, 0x1D, 0x1A, 0x5F, 0x09, 0x28,
	0x12, 0x26, 0x18, 0x58, 0x41, 0x0D, 0x70, 0x0E, 0x51, 0x5D, 0x0E, 0x18,
	0x27, 0x13, 0x5E, 0x5D, 0x0C, 0x5C, 0x18, 0x41, 0x1E, 0x7A, 0x0B, 0x2F,
	0x22, 0x52, 0x75, 0x2A, 0x33, 0x34, 0x1E, 0x7A, 0x03, 0x08, 0x56, 0x23,
	0x20, 0x0D, 0x15, 0x25, 0x5A, 0x03, 0x27, 0x59, 0x06, 0x59, 0x0A, 0x0F,
	0x59, 0x3A, 0x33, 0x2D, 0x1E, 0x53, 0x08, 0x02, 0x0C, 0x3A, 0x02, 0x03,
	0x40, 0x34, 0x54, 0x25, 0x0C, 0x0A, 0x17, 0x04, 0x08, 0x0A, 0x3F, 0x30,
	0x20, 0x14, 0x05, 0x5E, 0x33, 0x09, 0x14, 0x23, 0x21, 0x06, 0x09, 0x56,
	0x41, 0x2A, 0x17, 0x2B, 0x51, 0x21, 0x0E, 0x2F, 0x01, 0x31, 0x3E, 0x0A,
	0x73, 0x0F, 0x18, 0x18, 0x0F, 0x0A, 0x3C, 0x50, 0x2D, 0x3F, 0x28, 0x39,
	0x4A, 0x2D, 0x0A, 0x28, 0x20, 0x15, 0x38, 0x18, 0x04, 0x1B, 0x1B, 0x1F,
	0x5A, 0x77, 0x21, 0x16, 0x14, 0x05, 0x07, 0x25, 0x20, 0x1E, 0x3E, 0x09,
	0x16, 0x53, 0x5D, 0x32, 0x0A, 0x21, 0x10, 0x23, 0x1A, 0x0E, 0x0F, 0x56,
	0x3C, 0x3D, 0x38, 0x59, 0x29, 0x2C, 0x04, 0x34, 0x15, 0x0F, 0x18, 0x11,
	0x70, 0x03, 0x14, 0x1D, 0x23, 0x11, 0x59, 0x17, 0x59, 0x5E, 0x01, 0x24,
	0x13, 0x1D, 0x33, 0x73, 0x3B, 0x05, 0x2F, 0x12, 0x31, 0x5F, 0x52, 0x21,
	0x32, 0x13, 0x27, 0x00, 0x25, 0x27, 0x2E, 0x2D, 0x27, 0x14, 0x04, 0x74,
	0x1E, 0x05, 0x05, 0x21, 0x0D, 0x02, 0x0C, 0x3C, 0x18, 0x2E, 0x15, 0x06,
	0x0B, 0x5F, 0x17, 0x1A, 0x33, 0x57, 0x26, 0x35, 0x19, 0x02, 0x56, 0x07,
	0x24, 0x5A, 0x56, 0x20, 0x3F, 0x38, 0x06, 0x31, 0x58, 0x24, 0x72, 0x09,
	0x28, 0x1F, 0x5E, 0x21, 0x04, 0x2B, 0x0C, 0x29, 0x7A, 0x03, 0x0C, 0x56,
	0x3A, 0x12, 0x2F, 0x30, 0x2B, 0x38, 0x7B, 0x03, 0x06, 0x08, 0x39, 0x13,
	0x1A, 0x59, 0x5A, 0x1C, 0x2B, 0x00, 0x0F, 0x1B, 0x31, 0x0B, 0x2B, 0x05,
	0x16, 0x59, 0x2D, 0x1F, 0x31, 0x17, 0x11, 0x71, 0x09, 0x0B, 0x1D, 0x02,
	0x21, 0x1F, 0x09, 0x45, 0x1A, 0x29, 0x39, 0x12, 0x45, 0x5F, 0x36, 0x28,
	0x56, 0x00, 0x3D, 0x1B, 0x5E, 0x16, 0x1B, 0x3E, 0x0D, 0x3F, 0x25, 0x5C,
	0x3F, 0x74, 0x0F, 0x59, 0x0B, 0x2C, 0x05, 0x3E, 0x07, 0x5C, 0x38, 0x70,
	0x3B, 0x56, 0x5B, 0x01, 0x2F, 0x23, 0x22, 0x3B, 0x59, 0x75, 0x5C, 0x05,
	0x5D, 0x3A, 0x0E, 0x03, 0x39, 0x06, 0x59, 0x32, 0x35, 0x15, 0x39, 0x2F,
	0x09, 0x24, 0x50, 0x22, 0x0F, 0x2B, 0x1F, 0x04, 0x37, 0x0A, 0x23, 0x58,
	0x02, 0x0B, 0x39, 0x0B, 0x08, 0x51, 0x00, 0x5C, 0x06, 0x22, 0x4E, 0x27,
	0x32, 0x20, 0x0B, 0x52, 0x0D, 0x2A, 0x27, 0x54, 0x06, 0x0C, 0x2F, 0x31,
	0x0E, 0x2C, 0x39, 0x3F, 0x77, 0x2F, 0x56, 0x34, 0x24, 0x7A, 0x23, 0x39,
	0x08, 0x38, 0x07, 0x2B, 0x27, 0x59, 0x2F, 0x25, 0x07, 0x32, 0x23, 0x3D,
	0x16, 0x5F, 0x28, 0x2D, 0x52, 0x10, 0x34, 0x58, 0x5F, 0x26, 0x1B, 0x29,
	0x57, 0x18, 0x3B, 0x75, 0x1D, 0x34, 0x5E, 0x21, 0x73, 0x25, 0x3B, 0x45,
	0x5D, 0x32, 0x3D, 0x24, 0x0F, 0x19, 0x3A, 0x0E, 0x05, 0x14, 0x04, 0x07,
	0x06, 0x4E, 0x3F, 0x2C, 0x17, 0x1D, 0x0D, 0x07, 0x05, 0x34, 0x3A, 0x0D,
	0x24, 0x5C, 0x0C, 0x5A, 0x0E, 0x1A, 0x1E, 0x0F, 0x3C, 0x4A, 0x45, 0x33,
	0x3B, 0x14, 0x36, 0x3E, 0x3A, 0x25, 0x23, 0x39, 0x5D, 0x1C, 0x70, 0x06,
	0x2B, 0x2F, 0x5E, 0x14, 0x0E, 0x19, 0x2B, 0x2F, 0x3B, 0x28, 0x2C, 0x17,
	0x08, 0x07, 0x22, 0x35, 0x18, 0x00, 0x2A, 0x09, 0x0F, 0x1A, 0x31, 0x6D,
	0x25, 0x26, 0x25, 0x0C, 0x24, 0x1C, 0x2D, 0x36, 0x19, 0x37, 0x29, 0x15,
	0x09, 0x26, 0x25, 0x0A, 0x0E, 0x24, 0x21, 0x7A, 0x1D, 0x39, 0x5D, 0x21,
	0x6D, 0x20, 0x2F, 0x0F, 0x44, 0x33, 0x15, 0x07, 0x06, 0x1A, 0x06, 0x2A,
	0x10, 0x56, 0x5C, 0x1A, 0x2F, 0x57, 0x2D, 0x59, 0x70, 0x58, 0x29, 0x5F,
	0x3E, 0x0C, 0x2D, 0x56, 0x02, 0x29, 0x37, 0x38, 0x17, 0x3D, 0x5A, 0x08,
	0x39, 0x12, 0x05, 0x59, 0x7B, 0x09, 0x0B, 0x3E, 0x00, 0x05, 0x22, 0x06,
	0x1B, 0x24, 0x77, 0x19, 0x2F, 0x05, 0x12, 0x17, 0x2A, 0x24, 0x02, 0x2A,
	0x3A, 0x43, 0x4E, 0x17, 0x38, 0x1A, 0x39, 0x33, 0x3A, 0x26, 0x11, 0x00,
	0x0A, 0x1E, 0x31, 0x2F, 0x35, 0x16, 0x01, 0x22, 0x14, 0x58, 0x53, 0x0D,
	0x5D, 0x11, 0x19, 0x0C, 0x04, 0x44, 0x76, 0x07, 0x12, 0x29, 0x1D, 0x2E,
	0x39, 0x22, 0x58, 0x2A, 0x0B, 0x3C, 0x22, 0x05, 0x5D, 0x69, 0x20, 0x30,
	0x2A, 0x1A, 0x3A, 0x09, 0x58, 0x39, 0x08, 0x2F, 0x16, 0x04, 0x5F, 0x02,
	0x2E, 0x06, 0x31, 0x5D, 0x09, 0x25, 0x15, 0x37, 0x27, 0x26, 0x2D, 0x43,
	0x4E, 0x1D, 0x38, 0x07, 0x59, 0x29, 0x17, 0x53, 0x7B, 0x14, 0x14, 0x0B,
	0x53, 0x15, 0x39, 0x3B, 0x41, 0x1B, 0x2F, 0x2A, 0x0E, 0x0F, 0x3E, 0x11,
	0x1C, 0x24, 0x22, 0x06, 0x2C, 0x01, 0x28, 0x39, 0x00, 0x77, 0x06, 0x10,
	0x5F, 0x24, 0x0F, 0x07, 0x22, 0x17, 0x0D, 0x16, 0x35, 0x39, 0x2A, 0x5A,
	0x28, 0x3D, 0x0A, 0x01, 0x28, 0x35, 0x0A, 0x55, 0x5C, 0x40, 0x16, 0x5A,
	0x08, 0x5E, 0x44, 0x34, 0x20, 0x57, 0x29, 0x2E, 0x6D, 0x01, 0x2A, 0x03,
	0x3F, 0x36, 0x27, 0x05, 0x1A, 0x53, 0x69, 0x18, 0x35, 0x3E, 0x58, 0x13,
	0x38, 0x52, 0x5D, 0x00, 0x34, 0x2D, 0x0D, 0x24, 0x1E, 0x34, 0x54, 0x00,
	0x3E, 0x2C, 0x76, 0x3F, 0x0E, 0x37, 0x3B, 0x74, 0x34, 0x37, 0x5D, 0x3A,
	0x09, 0x0D, 0x56, 0x21, 0x12, 0x2F, 0x19, 0x0F, 0x41, 0x02, 0x0E, 0x26,
	0x36, 0x57, 0x33, 0x0B, 0x3C, 0x13, 0x5F, 0x11, 0x76, 0x28, 0x10, 0x38,
	0x5B, 0x70, 0x09, 0x35, 0x02, 0x29, 0x37, 0x3F, 0x29, 0x3E, 0x27, 0x2C,
	0x5D, 0x25, 0x45, 0x59, 0x1A, 0x25, 0x37, 0x2D, 0x09, 0x35, 0x47, 0x26,
	0x17, 0x18, 0x0A, 0x1D, 0x07, 0x39, 0x3D, 0x77, 0x21, 0x29, 0x0B, 0x06,
	0x71, 0x1A, 0x27, 0x26, 0x5D, 0x2A, 0x5F, 0x03, 0x1D, 0x33, 0x24, 0x5C,
	0x34, 0x1B, 0x40, 0x1B, 0x15, 0x12, 0x5A, 0x09, 0x13, 0x0A, 0x59, 0x5A,
	0x58, 0x69, 0x0A, 0x2C, 0x01, 0x1D, 0x76, 0x04, 0x54, 0x0B, 0x53, 0x31,
	0x3C, 0x55, 0x01, 0x20, 0x13, 0x20, 0x31, 0x16, 0x2A, 0x2D, 0x23, 0x34,
	0x5D, 0x12, 0x27, 0x19, 0x0C, 0x2B, 0x38, 0x3A, 0x3C, 0x11, 0x0C, 0x00,
	0x2D, 0x55, 0x11, 0x18, 0x04, 0x76, 0x02, 0x57, 0x2C, 0x0D, 0x15, 0x3C,
	0x52, 0x45, 0x29, 0x33, 0x47, 0x58, 0x58, 0x2E, 0x75, 0x01, 0x27, 0x00,
	0x44, 0x11, 0x21, 0x37, 0x45, 0x04, 0x27, 0x0B, 0x58, 0x5A, 0x52, 0x13,
	0x47, 0x36, 0x29, 0x05, 0x71, 0x29, 0x24, 0x0A, 0x13, 0x0A, 0x2A, 0x10,
	0x07, 0x5A, 0x2A, 0x3B, 0x36, 0x17, 0x29, 0x71, 0x54, 0x23, 0x5D, 0x00,
	0x24, 0x23, 0x06, 0x09, 0x3C, 0x14, 0x1B, 0x29, 0x25, 0x39, 0x6D, 0x3D,
	0x30, 0x3D, 0x5E, 0x2F, 0x38, 0x2B, 0x14, 0x07, 0x10, 0x24, 0x00, 0x0A,
	0x04, 0x71, 0x3C, 0x19, 0x45, 0x0D, 0x07, 0x09, 0x02, 0x09, 0x2C, 0x04,
	0x38, 0x58, 0x21, 0x31, 0x6D, 0x19, 0x2B, 0x5A, 0x2D, 0x7A, 0x00, 0x18,
	0x19, 0x29, 0x3A, 0x19, 0x1B, 0x39, 0x33, 0x7B, 0x55, 0x29, 0x01, 0x0D,
	0x37, 0x35, 0x25, 0x2D, 0x03, 0x6D, 0x0E, 0x35, 0x03, 0x13, 0x0E, 0x1C,
	0x04, 0x41, 0x1D, 0x2B, 0x55, 0x22, 0x03, 0x21, 0x7B, 0x2E, 0x50, 0x58,
	0x25, 0x75, 0x07, 0x38, 0x1B, 0x0C, 0x2C, 0x08, 0x25, 0x2F, 0x44, 0x26,
	0x26, 0x27, 0x5B, 0x3D, 0x71, 0x07, 0x59, 0x26, 0x19, 0x03, 0x54, 0x34,
	0x25, 0x26, 0x77, 0x0F, 0x57, 0x07, 0x20, 0x20, 0x1D, 0x02, 0x5D, 0x07,
	0x2F, 0x3E, 0x0A, 0x5E, 0x22, 0x3A, 0x2F, 0x05, 0x56, 0x00, 0x38, 0x1F,
	0x28, 0x14, 0x5D, 0x69, 0x06, 0x4A, 0x04, 0x52, 0x13, 0x5D, 0x28, 0x17,
	0x26, 0x6D, 0x54, 0x0E, 0x58, 0x2C, 0x37, 0x59, 0x13, 0x2B, 0x52, 0x31,
	0x08, 0x0C, 0x2F, 0x3D, 0x35, 0x43, 0x14, 0x0A, 0x52, 0x0C, 0x59, 0x51,
	0x59, 0x3B, 0x2E, 0x47, 0x58, 0x1C, 0x09, 0x25, 0x18, 0x0F, 0x45, 0x26,
	0x34, 0x3B, 0x52, 0x2F, 0x1D, 0x09, 0x43, 0x59, 0x05, 0x09, 0x05, 0x5F,
	0x2D, 0x0D, 0x5D, 0x7A, 0x07, 0x52, 0x28, 0x21, 0x74, 0x24, 0x0D, 0x2C,
	0x5A, 0x35, 0x0A, 0x59, 0x1E, 0x0C, 0x34, 0x43, 0x18, 0x20, 0x01, 0x75,
	0x0E, 0x17, 0x14, 0x01, 0x32, 0x3C, 0x50, 0x5D, 0x31, 0x05, 0x47, 0x2B,
	0x1D, 0x3F, 0x21, 0x1B, 0x14, 0x5D, 0x19, 0x1A, 0x39, 0x04, 0x22, 0x1F,
	0x7A, 0x0F, 0x0B, 0x0C, 0x2D, 0x2C, 0x3B, 0x0F, 0x28, 0x33, 0x2B, 0x5B,
	0x11, 0x1D, 0x31, 0x14, 0x0A, 0x4A, 0x36, 0x0F, 0x75, 0x15, 0x57, 0x59,
	0x0E, 0x7B, 0x3F, 0x25, 0x1A, 0x0E, 0x77, 0x07, 0x09, 0x59, 0x07, 0x03,
	0x0E, 0x08, 0x16, 0x28, 0x07, 0x47, 0x2B, 0x21, 0x02, 0x73, 0x18, 0x53,
	0x03, 0x20, 0x15, 0x2B, 0x07, 0x0B, 0x3B, 0x24, 0x1D, 0x0C, 0x5F, 0x09,
	0x2C, 0x1A, 0x18, 0x1A, 0x24, 0x3B, 0x47, 0x28, 0x58, 0x1D, 0x21, 0x5E,
	0x29, 0x22, 0x3D, 0x35, 0x07, 0x37, 0x06, 0x53, 0x1B, 0x15, 0x05, 0x1B,
	0x23, 0x31, 0x21, 0x51, 0x01, 0x2A, 0x71, 0x47, 0x56, 0x56, 0x29, 0x7B,
	0x3D, 0x59, 0x2D, 0x1F, 0x37, 0x27, 0x0C, 0x21, 0x3E, 0x38, 0x5B, 0x02,
	0x3A, 0x2C, 0x3A, 0x5F, 0x22, 0x58, 0x0C, 0x20, 0x3B, 0x08, 0x3F, 0x03,
	0x08, 0x23, 0x36, 0x5F, 0x13, 0x34, 0x5C, 0x0B, 0x41, 0x1F, 0x0E, 0x1A,
	0x26, 0x2D, 0x5C, 0x08, 0x5E, 0x57, 0x1D, 0x2F, 0x3B, 0x5C, 0x02, 0x1E,
	0x3E, 0x2A, 0x3E, 0x31, 0x17, 0x53, 0x37, 0x2A, 0x16, 0x16, 0x58, 0x29,
	0x00, 0x18, 0x5A, 0x25, 0x28, 0x0A, 0x10, 0x0D, 0x08, 0x37, 0x2E, 0x53,
	0x1A, 0x21, 0x27, 0x3D, 0x26, 0x03, 0x27, 0x77, 0x07, 0x11, 0x27, 0x27,
	0x38, 0x0D, 0x54, 0x5A, 0x3F, 0x2E, 0x15, 0x55, 0x26, 0x19, 0x69, 0x28,
	0x0D, 0x27, 0x52, 0x01, 0x15, 0x22, 0x59, 0x24, 0x35, 0x0A, 0x25, 0x3A,
	0x0E, 0x0C, 0x3B, 0x13, 0x29, 0x59, 0x7B, 0x26, 0x31, 0x01, 0x38, 0x30,
	0x5E, 0x34, 0x5E, 0x3A, 0x72, 0x0B, 0x30, 0x34, 0x59, 0x69, 0x1F, 0x0C,
	0x39, 0x1C, 0x6D, 0x21, 0x1B, 0x03, 0x5C, 0x23, 0x27, 0x50, 0x0D, 0x1F,
	0x10, 0x0F, 0x2B, 0x1B, 0x12, 0x09, 0x3B, 0x2D, 0x19, 0x0C, 0x09, 0x3D,
	0x2C, 0x0C, 0x0A, 0x0D, 0x16, 0x2D, 0x5A, 0x3B, 0x0D, 0x39, 0x0F, 0x27,
	0x1C, 0x2D, 0x28, 0x59, 0x0B, 0x19, 0x37, 0x2A, 0x54, 0x3D, 0x3B, 0x26,
	0x07, 0x27, 0x1A, 0x2D, 0x74, 0x0B, 0x2C, 0x17, 0x21, 0x71, 0x59, 0x2A,
	0x20, 0x09, 0x37, 0x2E, 0x4A, 0x00, 0x31, 0x70, 0x5F, 0x59, 0x59, 0x44,
	0x18, 0x43, 0x0D, 0x20, 0x04, 0x21, 0x00, 0x4A, 0x2F, 0x2F, 0x0E, 0x3E,
	0x0F, 0x5A, 0x26, 0x07, 0x29, 0x33, 0x36, 0x3B, 0x20, 0x5F, 0x28, 0x1D,
	0x1D, 0x38, 0x43, 0x24, 0x56, 0x59, 0x34, 0x59, 0x4E, 0x17, 0x24, 0x6D,
	0x14, 0x12, 0x3A, 0x53, 0x15, 0x1F, 0x56, 0x25, 0x27, 0x3B, 0x02, 0x55,
	0x2D, 0x0D, 0x26, 0x14, 0x2F, 0x36, 0x23, 0x71, 0x3E, 0x4E, 0x2B, 0x32,
	0x75, 0x09, 0x2C, 0x5C, 0x05, 0x17, 0x55, 0x57, 0x39, 0x02, 0x23, 0x09,
	0x31, 0x5F, 0x08, 0x0A, 0x34, 0x1B, 0x1E, 0x2A, 0x1A, 0x55, 0x37, 0x02,
	0x26, 0x2C, 0x39, 0x0A, 0x3E, 0x40, 0x2A, 0x2D, 0x2F, 0x45, 0x26, 0x2E,
	0x3F, 0x51, 0x56, 0x40, 0x3B, 0x43, 0x10, 0x29, 0x00, 0x75, 0x14, 0x58,
	0x3D, 0x3B, 0x75, 0x21, 0x58, 0x57, 0x0A, 0x38, 0x06, 0x0E, 0x20, 0x01,
	0x2A, 0x3C, 0x07, 0x34, 0x44, 0x29, 0x5B, 0x51, 0x3A, 0x1C, 0x30, 0x24,
	0x05, 0x3C, 0x58, 0x31, 0x04, 0x2E, 0x04, 0x2E, 0x3A, 0x3E, 0x31, 0x18,
	0x0F, 0x1A, 0x08, 0x0B, 0x00, 0x11, 0x16, 0x1E, 0x07, 0x0C, 0x20, 0x1B,
	0x08, 0x00, 0x05, 0x03, 0x2C, 0x35, 0x0D, 0x0A, 0x1A, 0x37, 0x25, 0x32,
	0x08, 0x19, 0x28, 0x3D, 0x59, 0x14, 0x1E, 0x09, 0x59, 0x07, 0x0A, 0x28,
	0x38, 0x23, 0x4A, 0x5F, 0x5F, 0x7A, 0x0B, 0x59, 0x59, 0x59, 0x32, 0x58,
	0x52, 0x18, 0x3A, 0x6D, 0x23, 0x2E, 0x3C, 0x08, 0x00, 0x0B, 0x24, 0x20,
	0x5D, 0x0A, 0x3A, 0x2E, 0x38, 0x3C, 0x27, 0x0A, 0x29, 0x0A, 0x40, 0x24,
	0x09, 0x30, 0x09, 0x0F, 0x2B, 0x07, 0x35, 0x26, 0x19, 0x18, 0x1C, 0x28,
	0x57, 0x5D, 0x1B, 0x1B, 0x07, 0x0A, 0x11, 0x11, 0x1B, 0x28, 0x59, 0x04,
	0x16, 0x14, 0x0E, 0x26, 0x12, 0x20, 0x14, 0x1B, 0x05, 0x3A, 0x04, 0x55,
	0x54, 0x08, 0x39, 0x0C, 0x14, 0x2E, 0x20, 0x3B, 0x0E, 0x0A, 0x29, 0x5F,
	0x04, 0x0C, 0x5C, 0x32, 0x21, 0x1F, 0x14, 0x0B, 0x2B, 0x58, 0x19, 0x17,
	0x0E, 0x18, 0x2C, 0x1B, 0x34, 0x2B, 0x05, 0x39, 0x0A, 0x08, 0x0D, 0x10,
	0x57, 0x11, 0x71, 0x09, 0x20, 0x0D, 0x1A, 0x31, 0x2E, 0x3B, 0x36, 0x31,
	0x27, 0x38, 0x36, 0x37, 0x3B, 0x69, 0x54, 0x0B, 0x5C, 0x3E, 0x2C, 0x00,
	0x24, 0x5A, 0x2D, 0x20, 0x5C, 0x10, 0x3D, 0x38, 0x08, 0x25, 0x07, 0x08,
	0x0A, 0x0A, 0x28, 0x55, 0x14, 0x38, 0x72, 0x23, 0x3B, 0x1A, 0x58, 0x20,
	0x58, 0x13, 0x2A, 0x3A, 0x20, 0x16, 0x23, 0x1D, 0x00, 0x26, 0x26, 0x25,
	0x2B, 0x00, 0x2D, 0x2A, 0x2F, 0x2C, 0x05, 0x07, 0x0F, 0x1B, 0x1C, 0x3B,
	0x13, 0x2D, 0x0D, 0x45, 0x01, 0x2D, 0x02, 0x31, 0x14, 0x13, 0x14, 0x5C,
	0x4A, 0x59, 0x0F, 0x0E, 0x19, 0x23, 0x22, 0x26, 0x76, 0x47, 0x52, 0x08,
	0x5B, 0x12, 0x3F, 0x4E, 0x27, 0x2C, 0x69, 0x0A, 0x10, 0x17, 0x3A, 0x25,
	0x15, 0x33, 0x45, 0x5C, 0x77, 0x29, 0x59, 0x1F, 0x23, 0x29, 0x5E, 0x2A,
	0x3A, 0x04, 0x15, 0x14, 0x25, 0x5C, 0x53, 0x0E, 0x5E, 0x30, 0x0B, 0x0C,
	0x20, 0x15, 0x13, 0x23, 0x1E, 0x32, 0x1F, 0x02, 0x27, 0x22, 0x11, 0x55,
	0x3B, 0x5F, 0x27, 0x04, 0x22, 0x07, 0x57, 0x20, 0x0C, 0x04, 0x08, 0x3B,
	0x0C, 0x2F, 0x5A, 0x0F, 0x08, 0x2E, 0x24, 0x19, 0x23, 0x22, 0x0D, 0x21,
	0x58, 0x37, 0x37, 0x12, 0x08, 0x58, 0x23, 0x17, 0x2C, 0x73, 0x3F, 0x35,
	0x57, 0x38, 0x36, 0x1E, 0x08, 0x1E, 0x38, 0x04, 0x14, 0x0B, 0x3A, 0x0A,
	0x6D, 0x19, 0x0F, 0x23, 0x02, 0x12, 0x01, 0x0B, 0x3F, 0x11, 0x74, 0x2A,
	0x0A, 0x36, 0x3D, 0x23, 0x1D, 0x12, 0x3E, 0x09, 0x6D, 0x35, 0x0B, 0x5A,
	0x5E, 0x06, 0x0B, 0x30, 0x09, 0x2F, 0x12, 0x55, 0x53, 0x34, 0x3E, 0x1B,
	0x00, 0x2C, 0x25, 0x28, 0x2A, 0x00, 0x2D, 0x3F, 0x38, 0x03, 0x03, 0x18,
	0x1D, 0x38, 0x01, 0x54, 0x1B, 0x29, 0x20, 0x2F, 0x43, 0x53, 0x01, 0x20,
	0x0F, 0x1E, 0x2A, 0x09, 0x1C, 0x75, 0x04, 0x34, 0x1A, 0x05, 0x04, 0x23,
	0x59, 0x05, 0x12, 0x6D, 0x1F, 0x05, 0x24, 0x5C, 0x05, 0x0B, 0x2D, 0x17,
	0x08, 0x03, 0x3A, 0x1B, 0x5A, 0x13, 0x09, 0x03, 0x0E, 0x34, 0x23, 0x12,
	0x09, 0x07, 0x1D, 0x0C, 0x76, 0x2B, 0x29, 0x0D, 0x1D, 0x34, 0x2A, 0x31,
	0x0B, 0x39, 0x0F, 0x2F, 0x23, 0x3F, 0x1A, 0x1B, 0x06, 0x4A, 0x1B, 0x04,
	0x6D, 0x0B, 0x16, 0x27, 0x1E, 0x0B, 0x03, 0x16, 0x58, 0x03, 0x1B, 0x1B,
	0x24, 0x28, 0x53, 0x0C, 0x2D, 0x05, 0x1D, 0x20, 0x3A, 0x25, 0x50, 0x3C,
	0x08, 0x27, 0x21, 0x4A, 0x25, 0x09, 0x28, 0x43, 0x00, 0x02, 0x0D, 0x35,
	0x5E, 0x18, 0x1D, 0x2A, 0x00, 0x19, 0x25, 0x41, 0x20, 0x11, 0x00, 0x55,
	0x56, 0x29, 0x2D, 0x1C, 0x04, 0x29, 0x2A, 0x7A, 0x3C, 0x2E, 0x45, 0x2F,
	0x6D, 0x47, 0x53, 0x1B, 0x32, 0x0A, 0x05, 0x2C, 0x02, 0x23, 0x75, 0x0F,
	0x27, 0x3A, 0x1C, 0x76, 0x5C, 0x09, 0x3B, 0x53, 0x21, 0x26, 0x55, 0x59,
	0x1D, 0x21, 0x0F, 0x37, 0x59, 0x2F, 0x00, 0x20, 0x57, 0x36, 0x1D, 0x21,
	0x5A, 0x34, 0x28, 0x33, 0x69, 0x07, 0x05, 0x28, 0x5D, 0x11, 0x0A, 0x05,
	0x56, 0x03, 0x74, 0x54, 0x0F, 0x3B, 0x5C, 0x27, 0x06, 0x07, 0x0D, 0x3C,
	0x76, 0x2F, 0x54, 0x25, 0x18, 0x0A, 0x22, 0x59, 0x3B, 0x0D, 0x32, 0x09,
	0x57, 0x28, 0x5B, 0x70, 0x1A, 0x23, 0x27, 0x38, 0x12, 0x5F, 0x27, 0x5E,
	0x08, 0x2C, 0x2E, 0x4E, 0x29, 0x05, 0x76, 0x2E, 0x2B, 0x3E, 0x05, 0x35,
	0x08, 0x2D, 0x3D, 0x13, 0x0F, 0x06, 0x15, 0x57, 0x0F, 0x74, 0x38, 0x53,
	0x3F, 0x0A, 0x28, 0x38, 0x2F, 0x17, 0x18, 0x73, 0x5A, 0x0A, 0x19, 0x3B,
	0x37, 0x04, 0x37, 0x59, 0x28, 0x31, 0x28, 0x51, 0x5A, 0x5C, 0x0B, 0x5B,
	0x15, 0x38, 0x0F, 0x11, 0x2F, 0x15, 0x20, 0x08, 0x69, 0x3E, 0x4A, 0x25,
	0x5A, 0x27, 0x43, 0x50, 0x01, 0x33, 0x29, 0x22, 0x0C, 0x03, 0x29, 0x0C,
	0x0F, 0x27, 0x1C, 0x58, 0x0D, 0x59, 0x36, 0x0C, 0x5B, 0x74, 0x35, 0x11,
	0x59, 0x05, 0x0A, 0x08, 0x50, 0x04, 0x31, 0x21, 0x0D, 0x50, 0x5D, 0x3F,
	0x2A, 0x28, 0x37, 0x0B, 0x5B, 0x37, 0x0B, 0x2F, 0x24, 0x2E, 0x0C, 0x28,
	0x17, 0x3E, 0x13, 0x2C, 0x3C, 0x31, 0x59, 0x59, 0x23, 0x36, 0x24, 0x3F,
	0x07, 0x32, 0x59, 0x50, 0x2D, 0x07, 0x31, 0x5B, 0x51, 0x5C, 0x3B, 0x73,
	0x5F, 0x16, 0x01, 0x07, 0x7B, 0x05, 0x33, 0x59, 0x0E, 0x74, 0x24, 0x59,
	0x0C, 0x1A, 0x35, 0x0B, 0x30, 0x28, 0x29, 0x2E, 0x5E, 0x03, 0x57, 0x58,
	0x17, 0x22, 0x23, 0x0F, 0x1A, 0x0C, 0x34, 0x11, 0x41, 0x1B, 0x05, 0x43,
	0x19, 0x5C, 0x28, 0x00, 0x2E, 0x35, 0x5F, 0x24, 0x13, 0x3E, 0x0A, 0x37,
	0x31, 0x05, 0x35, 0x09, 0x57, 0x5A, 0x0C, 0x1E, 0x3B, 0x3E, 0x53, 0x69,
	0x19, 0x25, 0x56, 0x5C, 0x27, 0x2B, 0x22, 0x27, 0x12, 0x3A, 0x1F, 0x16,
	0x38, 0x1E, 0x76, 0x5F, 0x26, 0x2D, 0x21, 0x2B, 0x59, 0x30, 0x28, 0x2F,
	0x76, 0x24, 0x11, 0x2A, 0x18, 0x01, 0x3C, 0x2F, 0x2B, 0x0E, 0x35, 0x35,
	0x0A, 0x0C, 0x5C, 0x0A, 0x01, 0x05, 0x59, 0x06, 0x29, 0x20, 0x04, 0x00,
	0x09, 0x35, 0x55, 0x10, 0x19, 0x13, 0x73, 0x3D, 0x19, 0x23, 0x04, 0x0D,
	0x3D, 0x54, 0x3D, 0x40, 0x73, 0x47, 0x54, 0x23, 0x09, 0x35, 0x09, 0x08,
	0x57, 0x24, 0x70, 0x0B, 0x34, 0x3D, 0x09, 0x0E, 0x1F, 0x50, 0x22, 0x3B,
	0x3B, 0x25, 0x04, 0x0D, 0x5A, 0x29, 0x36, 0x17, 0x0C, 0x5C, 0x0E, 0x58,
	0x54, 0x28, 0x11, 0x21, 0x18, 0x03, 0x0C, 0x1E, 0x2A, 0x1C, 0x26, 0x58,
	0x52, 0x23, 0x15, 0x33, 0x03, 0x06, 0x20, 0x06, 0x12, 0x5C, 0x06, 0x34,
	0x2A, 0x0A, 0x08, 0x24, 0x15, 0x35, 0x1B, 0x41, 0x59, 0x15, 0x58, 0x23,
	0x41, 0x01, 0x31, 0x1C, 0x55, 0x3C, 0x13, 0x7B, 0x54, 0x23, 0x57, 0x04,
	0x0E, 0x19, 0x54, 0x24, 0x3F, 0x14, 0x2D, 0x4A, 0x26, 0x5D, 0x6D, 0x2A,
	0x00, 0x3A, 0x3C, 0x09, 0x29, 0x27, 0x5C, 0x06, 0x06, 0x3C, 0x0A, 0x2A,
	0x3C, 0x71, 0x08, 0x20, 0x20, 0x33, 0x14, 0x36, 0x0B, 0x26, 0x22, 0x69,
	0x5A, 0x00, 0x0A, 0x2A, 0x12, 0x1E, 0x14, 0x39, 0x1B, 0x37, 0x1A, 0x38,
	0x3A, 0x58, 0x7B, 0x02, 0x38, 0x21, 0x52, 0x09, 0x25, 0x37, 0x22, 0x1D,
	0x17, 0x5E, 0x18, 0x1B, 0x3F, 0x32, 0x22, 0x1B, 0x18, 0x59, 0x2E, 0x21,
	0x2D, 0x37, 0x24, 0x2D, 0x08, 0x10, 0x18, 0x07, 0x15, 0x1D, 0x2B, 0x0B,
	0x0E, 0x34, 0x5A, 0x38, 0x5C, 0x20, 0x0E, 0x28, 0x4E, 0x5B, 0x19, 0x26,
	0x23, 0x58, 0x0F, 0x0F, 0x2C, 0x08, 0x52, 0x3F, 0x02, 0x76, 0x25, 0x23,
	0x1E, 0x18, 0x76, 0x1F, 0x15, 0x5F, 0x1B, 0x10, 0x0A, 0x22, 0x36, 0x02,
	0x24, 0x5C, 0x50, 0x23, 0x3B, 0x07, 0x08, 0x08, 0x5D, 0x03, 0x27, 0x14,
	0x56, 0x22, 0x25, 0x2B, 0x1D, 0x34, 0x39, 0x39, 0x25, 0x5B, 0x32, 0x56,
	0x3A, 0x03, 0x29, 0x0E, 0x20, 0x1E, 0x28, 0x2B, 0x56, 0x1C, 0x52, 0x0F,
	0x47, 0x35, 0x57, 0x3B, 0x2C, 0x36, 0x53, 0x17, 0x2D, 0x20, 0x22, 0x54,
	0x3C, 0x12, 0x38, 0x04, 0x17, 0x41, 0x09, 0x7B, 0x5D, 0x55, 0x00, 0x25,
	0x12, 0x5C, 0x05, 0x07, 0x05, 0x6D, 0x47, 0x3B, 0x02, 0x07, 0x20, 0x5C,
	0x19, 0x29, 0x5C, 0x30, 0x5A, 0x4E, 0x0A, 0x23, 0x14, 0x06, 0x58, 0x41,
	0x2A, 0x2E, 0x58, 0x25, 0x29, 0x39, 0x0C, 0x3F, 0x57, 0x18, 0x32, 0x20,
	0x39, 0x27, 0x3C, 0x1E, 0x07, 0x0D, 0x50, 0x18, 0x5E, 0x18, 0x1E, 0x09,
	0x04, 0x3C, 0x28, 0x08, 0x0F, 0x29, 0x1E, 0x00, 0x34, 0x57, 0x0A, 0x04,
	0x30, 0x0F, 0x10, 0x5F, 0x18, 0x1B, 0x0A, 0x37, 0x1B, 0x33, 0x20, 0x5E,
	0x12, 0x2D, 0x5C, 0x1A, 0x21, 0x16, 0x2B, 0x1D, 0x2B, 0x1F, 0x2A, 0x28,
	0x09, 0x77, 0x0B, 0x27, 0x5F, 0x2A, 0x05, 0x3D, 0x23, 0x28, 0x28, 0x17,
	0x3C, 0x0F, 0x0C, 0x01, 0x34, 0x18, 0x51, 0x2B, 0x2D, 0x0F, 0x23, 0x07,
	0x1B, 0x1F, 0x2A, 0x59, 0x20, 0x0D, 0x02, 0x2E, 0x3B, 0x36, 0x2D, 0x5E,
	0x08, 0x20, 0x51, 0x1D, 0x52, 0x2F, 0x2F, 0x31, 0x3E, 0x3E, 0x38, 0x2B,
	0x23, 0x14, 0x52, 0x7A, 0x2D, 0x54, 0x5E, 0x1A, 0x30, 0x3F, 0x2F, 0x07,
	0x06, 0x0B, 0x08, 0x0D, 0x5A, 0x11, 0x23, 0x38, 0x07, 0x5D, 0x5B, 0x37,
	0x5F, 0x0C, 0x5C, 0x3B, 0x27, 0x5C, 0x58, 0x2F, 0x26, 0x08, 0x02, 0x2E,
	0x1A, 0x09, 0x77, 0x2A, 0x09, 0x5A, 0x07, 0x35, 0x1C, 0x16, 0x27, 0x1D,
	0x71, 0x0A, 0x2C, 0x27, 0x1E, 0x33, 0x5B, 0x0E, 0x59, 0x31, 0x71, 0x5C,
	0x51, 0x27, 0x3C, 0x11, 0x21, 0x13, 0x3B, 0x3C, 0x0D, 0x1C, 0x0E, 0x0D,
	0x00, 0x29, 0x1D, 0x2C, 0x1F, 0x12, 0x11, 0x04, 0x2E, 0x16, 0x1A, 0x0D,
	0x1E, 0x19, 0x0B, 0x5D, 0x77, 0x38, 0x2C, 0x09, 0x0A, 0x21, 0x00, 0x38,
	0x5D, 0x52, 0x37, 0x34, 0x2A, 0x04, 0x5F, 0x16, 0x0F, 0x2E, 0x3B, 0x0D,
	0x07, 0x55, 0x02, 0x5C, 0x01, 0x25, 0x59, 0x37, 0x2C, 0x08, 0x33, 0x15,
	0x00, 0x08, 0x58, 0x3B, 0x05, 0x2E, 0x2F, 0x52, 0x01, 0x18, 0x2D, 0x09,
	0x59, 0x04, 0x25, 0x35, 0x2B, 0x2F, 0x3A, 0x5C, 0x1B, 0x2D, 0x3D, 0x30,
	0x3E, 0x05, 0x37, 0x0E, 0x33, 0x3F, 0x36, 0x2F, 0x3E, 0x27, 0x38, 0x0B,
	0x23, 0x18, 0x31, 0x3F, 0x36, 0x37, 0x06, 0x3A, 0x20, 0x24, 0x06, 0x0F,
	0x0B, 0x0A, 0x07, 0x01, 0x26, 0x0A, 0x25, 0x10, 0x5B, 0x03, 0x05, 0x3C,
	0x59, 0x56, 0x03, 0x74, 0x25, 0x32, 0x2C, 0x1D, 0x0F, 0x1F, 0x12, 0x1B,
	0x5C, 0x28, 0x0E, 0x38, 0x05, 0x26, 0x16, 0x28, 0x0B, 0x03, 0x3F, 0x77,
	0x1A, 0x10, 0x2D, 0x01, 0x18, 0x24, 0x17, 0x57, 0x2C, 0x71, 0x25, 0x0F,
	0x5A, 0x24, 0x34, 0x5A, 0x15, 0x5B, 0x53, 0x36, 0x09, 0x04, 0x0B, 0x1D,
	0x2F, 0x14, 0x56, 0x29, 0x24, 0x71, 0x0D, 0x2F, 0x3B, 0x07, 0x27, 0x24,
	0x4A, 0x3E, 0x0A, 0x0A, 0x1B, 0x32, 0x20, 0x06, 0x33, 0x09, 0x53, 0x3F,
	0x1F, 0x09, 0x2F, 0x19, 0x22, 0x04, 0x26, 0x25, 0x2B, 0x39, 0x18, 0x28,
	0x34, 0x32, 0x3F, 0x44, 0x2B, 0x23, 0x03, 0x5F, 0x33, 0x72, 0x02, 0x04,
	0x5D, 0x07, 0x10, 0x14, 0x54, 0x39, 0x00, 0x2A, 0x59, 0x06, 0x41, 0x0F,
	0x30, 0x3F, 0x1B, 0x1E, 0x39, 0x34, 0x18, 0x37, 0x07, 0x12, 0x36, 0x58,
	0x2F, 0x2C, 0x05, 0x12, 0x20, 0x05, 0x1C, 0x08, 0x35, 0x23, 0x2D, 0x04,
	0x09, 0x73, 0x20, 0x14, 0x3E, 0x1B, 0x07, 0x01, 0x0E, 0x5A, 0x0E, 0x72,
	0x5E, 0x29, 0x1F, 0x23, 0x37, 0x28, 0x24, 0x24, 0x39, 0x0F, 0x3D, 0x0B,
	0x2F, 0x1F, 0x76, 0x05, 0x20, 0x19, 0x52, 0x0E, 0x09, 0x08, 0x26, 0x00,
	0x29, 0x08, 0x2C, 0x2D, 0x38, 0x33, 0x5C, 0x0D, 0x3E, 0x53, 0x01, 0x0A,
	0x2E, 0x39, 0x08, 0x21, 0x3D, 0x06, 0x1B, 0x53, 0x2F, 0x22, 0x38, 0x26,
	0x04, 0x06, 0x2E, 0x00, 0x27, 0x3B, 0x13, 0x59, 0x09, 0x39, 0x5D, 0x2C,
	0x5C, 0x2E, 0x3B, 0x3E, 0x0B, 0x07, 0x2A, 0x08, 0x5B, 0x01, 0x5E, 0x02,
	0x28, 0x28, 0x0B, 0x23, 0x38, 0x0C, 0x0E, 0x35, 0x5E, 0x18, 0x05, 0x2E,
	0x2C, 0x39, 0x2B, 0x2F, 0x0A, 0x00, 0x3B, 0x53, 0x28, 0x1E, 0x14, 0x5F,
	0x0D, 0x22, 0x40, 0x09, 0x20, 0x12, 0x25, 0x0C, 0x08, 0x3F, 0x20, 0x2A,
	0x09, 0x28, 0x55, 0x59, 0x26, 0x2E, 0x73, 0x2B, 0x11, 0x17, 0x05, 0x05,
	0x5B, 0x58, 0x21, 0x32, 0x7B, 0x00, 0x2C, 0x05, 0x0F, 0x7A, 0x2F, 0x2C,
	0x0F, 0x0E, 0x29, 0x25, 0x26, 0x2F, 0x44, 0x2A, 0x47, 0x4E, 0x2C, 0x1B,
	0x13, 0x3D, 0x09, 0x21, 0x3D, 0x76, 0x14, 0x0C, 0x1E, 0x11, 0x17, 0x1F,
	0x07, 0x2F, 0x03, 0x34, 0x00, 0x10, 0x06, 0x12, 0x74, 0x5F, 0x12, 0x3E,
	0x3D, 0x09, 0x3E, 0x36, 0x3D, 0x24, 0x0B, 0x0E, 0x1B, 0x0F, 0x29, 0x05,
	0x34, 0x03, 0x05, 0x0C, 0x21, 0x2E, 0x19, 0x05, 0x06, 0x16, 0x39, 0x0E,
	0x1F, 0x5A, 0x38, 0x25, 0x37, 0x1E, 0x0D, 0x73, 0x1F, 0x51, 0x5F, 0x32,
	0x08, 0x3B, 0x2B, 0x5F, 0x24, 0x28, 0x3E, 0x28, 0x56, 0x29, 0x37, 0x16,
	0x55, 0x1D, 0x1C, 0x72, 0x3D, 0x2C, 0x5F, 0x24, 0x2D, 0x26, 0x0E, 0x1A,
	0x1D, 0x6D, 0x04, 0x00, 0x0A, 0x05, 0x36, 0x06, 0x4A, 0x36, 0x21, 0x29,
	0x2F, 0x53, 0x3C, 0x29, 0x26, 0x43, 0x2B, 0x19, 0x09, 0x20, 0x3B, 0x09,
	0x41, 0x11, 0x77, 0x22, 0x27, 0x07, 0x04, 0x08, 0x47, 0x58, 0x17, 0x28,
	0x05, 0x5B, 0x14, 0x29, 0x2C, 0x73, 0x0A, 0x4A, 0x26, 0x18, 0x17, 0x02,
	0x0C, 0x5F, 0x1D, 0x76, 0x39, 0x11, 0x24, 0x1F, 0x26, 0x21, 0x55, 0x19,
	0x5C, 0x34, 0x08, 0x4A, 0x1C, 0x44, 0x33, 0x34, 0x0C, 0x5B, 0x07, 0x30,
	0x02, 0x30, 0x02, 0x38, 0x7A, 0x01, 0x03, 0x29, 0x5F, 0x29, 0x1E, 0x53,
	0x0D, 0x25, 0x13, 0x07, 0x32, 0x20, 0x02, 0x2A, 0x03, 0x1B, 0x1B, 0x33,
	0x0A, 0x24, 0x39, 0x24, 0x21, 0x72, 0x38, 0x17, 0x0A, 0x3A, 0x2E, 0x47,
	0x2A, 0x14, 0x2D, 0x26, 0x55, 0x34, 0x0F, 0x3B, 0x07, 0x3C, 0x59, 0x07,
	0x18, 0x04, 0x5E, 0x02, 0x56, 0x0D, 0x05, 0x5C, 0x29, 0x3C, 0x5C, 0x36,
	0x29, 0x59, 0x08, 0x19, 0x2C, 0x3B, 0x19, 0x56, 0x19, 0x08, 0x23, 0x2F,
	0x04, 0x58, 0x15, 0x15, 0x59, 0x0C, 0x2D, 0x0D, 0x22, 0x11, 0x5B, 0x5A,
	0x0F, 0x04, 0x25, 0x34, 0x59, 0x04, 0x29, 0x29, 0x07, 0x24, 0x35, 0x05,
	0x4A, 0x3C, 0x24, 0x17, 0x22, 0x20, 0x26, 0x1F, 0x00, 0x36, 0x30, 0x58,
	0x04, 0x0B, 0x0A, 0x2B, 0x1B, 0x13, 0x38, 0x15, 0x2D, 0x00, 0x3A, 0x35,
	0x2D, 0x56, 0x5F, 0x1F, 0x37, 0x22, 0x56, 0x0C, 0x3C, 0x2E, 0x06, 0x05,
	0x2D, 0x24, 0x38, 0x3E, 0x0E, 0x04, 0x53, 0x01, 0x18, 0x00, 0x3B, 0x22,
	0x15, 0x22, 0x58, 0x59, 0x20, 0x14, 0x5C, 0x57, 0x1A, 0x0D, 0x04, 0x54,
	0x0D, 0x14, 0x21, 0x16, 0x0F, 0x2B, 0x2F, 0x3C, 0x0B, 0x5A, 0x4A, 0x04,
	0x1E, 0x05, 0x58, 0x51, 0x20, 0x5E, 0x2D, 0x14, 0x08, 0x2A, 0x04, 0x28,
	0x35, 0x0A, 0x03, 0x31, 0x0E, 0x58, 0x06, 0x0C, 0x08, 0x24, 0x3F, 0x23,
	0x5C, 0x03, 0x74, 0x26, 0x18, 0x37, 0x3F, 0x35, 0x1D, 0x2E, 0x25, 0x28,
	0x13, 0x20, 0x37, 0x5B, 0x3C, 0x2A, 0x1C, 0x59, 0x28, 0x19, 0x14, 0x0A,
	0x09, 0x59, 0x33, 0x18, 0x5C, 0x39, 0x0C, 0x3E, 0x0B, 0x38, 0x30, 0x59,
	0x0C, 0x29, 0x09, 0x2F, 0x3A, 0x01, 0x29, 0x3F, 0x25, 0x24, 0x1E, 0x21,
	0x5D, 0x0E, 0x07, 0x5A, 0x07, 0x3A, 0x57, 0x36, 0x01, 0x77, 0x38, 0x0E,
	0x1E, 0x28, 0x27, 0x1D, 0x34, 0x57, 0x21, 0x1B, 0x00, 0x0B, 0x5F, 0x5B,
	0x7B, 0x3F, 0x37, 0x39, 0x1F, 0x13, 0x5F, 0x23, 0x09, 0x59, 0x34, 0x24,
	0x53, 0x21, 0x3D, 0x2D, 0x58, 0x15, 0x01, 0x2A, 0x7B, 0x39, 0x17, 0x01,
	0x00, 0x26, 0x03, 0x11, 0x3E, 0x24, 0x70, 0x2B, 0x2E, 0x07, 0x03, 0x72,
	0x3B, 0x13, 0x14, 0x5B, 0x2F, 0x0B, 0x38, 0x2F, 0x1F, 0x01, 0x16, 0x4A,
	0x05, 0x5E, 0x2C, 0x3B, 0x23, 0x57, 0x11, 0x09, 0x0E, 0x20, 0x28, 0x1D,
	0x2F, 0x1E, 0x2A, 0x1F, 0x2E, 0x2A, 0x1D, 0x51, 0x1C, 0x33, 0x2C, 0x2B,
	0x0E, 0x21, 0x44, 0x30, 0x19, 0x36, 0x29, 0x2E, 0x35, 0x59, 0x52, 0x3B,
	0x25, 0x26, 0x47, 0x2C, 0x09, 0x29, 0x2E, 0x55, 0x52, 0x17, 0x03, 0x3A,
	0x59, 0x36, 0x0B, 0x31, 0x2F, 0x2A, 0x32, 0x37, 0x1D, 0x08, 0x3B, 0x2B,
	0x59, 0x5D, 0x7B, 0x16, 0x2D, 0x01, 0x24, 0x29, 0x1D, 0x58, 0x1A, 0x2D,
	0x2C, 0x16, 0x2C, 0x0C, 0x12, 0x2A, 0x1F, 0x2A, 0x0A, 0x1A, 0x24, 0x20,
	0x30, 0x0D, 0x02, 0x28, 0x18, 0x05, 0x03, 0x5A, 0x7A, 0x43, 0x22, 0x1E,
	0x31, 0x29, 0x2B, 0x12, 0x0C, 0x01, 0x17, 0x02, 0x51, 0x02, 0x08, 0x3A,
	0x47, 0x0E, 0x2A, 0x04, 0x29, 0x5B, 0x2B, 0x1E, 0x1F, 0x37, 0x3F, 0x20,
	0x29, 0x2E, 0x74, 0x25, 0x55, 0x06, 0x1D, 0x2F, 0x36, 0x29, 0x29, 0x59,
	0x13, 0x26, 0x19, 0x2C, 0x2D, 0x7A, 0x25, 0x56, 0x5D, 0x58, 0x16, 0x21,
	0x0A, 0x1D, 0x1D, 0x20, 0x00, 0x23, 0x3A, 0x27, 0x73, 0x1C, 0x2C, 0x22,
	0x38, 0x0C, 0x35, 0x2C, 0x2B, 0x3D, 0x21, 0x3A, 0x0B, 0x0F, 0x2A, 0x2B,
	0x2F, 0x4A, 0x25, 0x3F, 0x34, 0x14, 0x08, 0x2C, 0x12, 0x26, 0x47, 0x23,
	0x24, 0x39, 0x34, 0x58, 0x25, 0x3A, 0x06, 0x0B, 0x34, 0x19, 0x03, 0x24,
	0x37, 0x3B, 0x0E, 0x23, 0x52, 0x33, 0x36, 0x56, 0x2A, 0x1C, 0x2C, 0x59,
	0x2B, 0x56, 0x3A, 0x14, 0x00, 0x57, 0x3E, 0x1F, 0x32, 0x1D, 0x19, 0x1F,
	0x58, 0x77, 0x06, 0x08, 0x45, 0x11, 0x3B, 0x14, 0x04, 0x1E, 0x2C, 0x12,
	0x08, 0x50, 0x58, 0x2E, 0x27, 0x1E, 0x2A, 0x5A, 0x18, 0x13, 0x28, 0x32,
	0x5D, 0x02, 0x33, 0x2D, 0x38, 0x3E, 0x22, 0x05, 0x5C, 0x50, 0x14, 0x1B,
	0x15, 0x43, 0x23, 0x29, 0x52, 0x04, 0x3B, 0x35, 0x5E, 0x5C, 0x03, 0x08,
	0x0B, 0x17, 0x11, 0x18, 0x5B, 0x55, 0x0F, 0x0E, 0x74, 0x3D, 0x27, 0x3C,
	0x21, 0x2C, 0x55, 0x24, 0x0A, 0x00, 0x0B, 0x0B, 0x51, 0x37, 0x1A, 0x31,
	0x23, 0x59, 0x05, 0x1E, 0x2F, 0x58, 0x0D, 0x02, 0x3B, 0x12, 0x07, 0x07,
	0x5F, 0x08, 0x76, 0x5B, 0x35, 0x3B, 0x32, 0x0D, 0x58, 0x55, 0x18, 0x1C,
	0x12, 0x2F, 0x06, 0x03, 0x3B, 0x23, 0x20, 0x0C, 0x1C, 0x23, 0x16, 0x16,
	0x53, 0x5E, 0x3F, 0x34, 0x5C, 0x27, 0x3D, 0x3C, 0x20, 0x2D, 0x04, 0x02,
	0x28, 0x01, 0x02, 0x37, 0x36, 0x53, 0x03, 0x3F, 0x56, 0x0F, 0x12, 0x28,
	0x1D, 0x2F, 0x5D, 0x2E, 0x0D, 0x5B, 0x04, 0x24, 0x08, 0x23, 0x0D, 0x33,
	0x04, 0x5D, 0x0F, 0x5F, 0x18, 0x1E, 0x5A, 0x2A, 0x05, 0x23, 0x56, 0x1D,
	0x7A, 0x08, 0x17, 0x1C, 0x05, 0x0F, 0x3C, 0x2F, 0x39, 0x3B, 0x08, 0x2B,
	0x10, 0x1E, 0x1C, 0x3A, 0x1D, 0x30, 0x20, 0x19, 0x0A, 0x22, 0x4E, 0x24,
	0x01, 0x14, 0x0B, 0x03, 0x2A, 0x5E, 0x7B, 0x02, 0x2C, 0x2B, 0x29, 0x7B,
	0x3D, 0x56, 0x3B, 0x19, 0x7B, 0x05, 0x06, 0x58, 0x1D, 0x16, 0x0D, 0x0D,
	0x3B, 0x05, 0x14, 0x5C, 0x31, 0x01, 0x0D, 0x69, 0x1E, 0x09, 0x21, 0x11,
	0x27, 0x47, 0x26, 0x56, 0x08, 0x69, 0x0A, 0x39, 0x23, 0x5F, 0x28, 0x3C,
	0x56, 0x5A, 0x3E, 0x31, 0x1A, 0x58, 0x01, 0x31, 0x21, 0x0B, 0x08, 0x27,
	0x3A, 0x35, 0x26, 0x24, 0x26, 0x1C, 0x71, 0x1C, 0x0F, 0x3C, 0x3D, 0x24,
	0x0E, 0x17, 0x39, 0x2C, 0x17, 0x43, 0x29, 0x2B, 0x5F, 0x2D, 0x35, 0x2C,
	0x02, 0x18, 0x25, 0x34, 0x13, 0x2C, 0x04, 0x36, 0x09, 0x06, 0x1C, 0x1D,
	0x3A, 0x2A, 0x31, 0x27, 0x28, 0x70, 0x1B, 0x00, 0x37, 0x53, 0x03, 0x0E,
	0x38, 0x25, 0x03, 0x27, 0x5E, 0x30, 0x07, 0x06, 0x34, 0x08, 0x28, 0x3A,
	0x0E, 0x75, 0x5D, 0x11, 0x22, 0x27, 0x76, 0x21, 0x51, 0x20, 0x28, 0x06,
	0x3F, 0x35, 0x2F, 0x28, 0x0A, 0x2A, 0x15, 0x19, 0x12, 0x15, 0x1F, 0x19,
	0x21, 0x1E, 0x0C, 0x58, 0x0C, 0x06, 0x2D, 0x06, 0x3D, 0x13, 0x02, 0x18,
	0x2C, 0x07, 0x25, 0x2B, 0x05, 0x24, 0x47, 0x2E, 0x1E, 0x11, 0x7A, 0x23,
	0x06, 0x02, 0x05, 0x1B, 0x05, 0x4E, 0x29, 0x24, 0x29, 0x34, 0x58, 0x2B,
	0x52, 0x07, 0x59, 0x2E, 0x5E, 0x3F, 0x2F, 0x0A, 0x13, 0x27, 0x44, 0x21,
	0x54, 0x0B, 0x26, 0x08, 0x2A, 0x0E, 0x02, 0x0B, 0x08, 0x7B, 0x23, 0x28,
	0x0C, 0x5B, 0x1A, 0x5F, 0x0D, 0x34, 0x22, 0x76, 0x29, 0x57, 0x37, 0x39,
	0x07, 0x0A, 0x52, 0x24, 0x21, 0x1A, 0x08, 0x2D, 0x19, 0x03, 0x2F, 0x24,
	0x15, 0x3B, 0x53, 0x73, 0x19, 0x0A, 0x28, 0x28, 0x01, 0x35, 0x58, 0x2D,
	0x21, 0x09, 0x06, 0x2B, 0x5C, 0x33, 0x11, 0x1C, 0x16, 0x00, 0x08, 0x35,
	0x36, 0x35, 0x5F, 0x3D, 0x2E, 0x35, 0x17, 0x1B, 0x22, 0x35, 0x3F, 0x19,
	0x0F, 0x1D, 0x08, 0x0B, 0x29, 0x27, 0x28, 0x00, 0x09, 0x57, 0x2F, 0x25,
	0x7B, 0x5A, 0x05, 0x2D, 0x58, 0x27, 0x3A, 0x4E, 0x24, 0x23, 0x30, 0x34,
	0x30, 0x58, 0x29, 0x7A, 0x34, 0x25, 0x18, 0x38, 0x34, 0x5F, 0x55, 0x0F,
	0x11, 0x69, 0x27, 0x0D, 0x1D, 0x38, 0x3A, 0x1D, 0x31, 0x37, 0x07, 0x73,
	0x23, 0x50, 0x0F, 0x05, 0x11, 0x5A, 0x09, 0x08, 0x1A, 0x04, 0x16, 0x27,
	0x05, 0x0E, 0x20, 0x18, 0x35, 0x06, 0x3D, 0x1A, 0x43, 0x30, 0x18, 0x3F,
	0x01, 0x5E, 0x2D, 0x1A, 0x0D, 0x31, 0x3A, 0x10, 0x5F, 0x5D, 0x30, 0x34,
	0x56, 0x02, 0x1C, 0x74, 0x22, 0x15, 0x1D, 0x25, 0x23, 0x3E, 0x23, 0x22,
	0x1F, 0x15, 0x3E, 0x06, 0x2D, 0x06, 0x20, 0x07, 0x2A, 0x18, 0x59, 0x15,
	0x34, 0x15, 0x14, 0x13, 0x06, 0x58, 0x03, 0x3A, 0x5B, 0x29, 0x22, 0x18,
	0x2A, 0x3B, 0x21, 0x00, 0x08, 0x58, 0x1D, 0x35, 0x5E, 0x20, 0x01, 0x1E,
	0x25, 0x1E, 0x59, 0x5B, 0x28, 0x12, 0x1F, 0x4E, 0x08, 0x2C, 0x03, 0x05,
	0x58, 0x1F, 0x01, 0x28, 0x02, 0x39, 0x45, 0x1A, 0x2B, 0x0A, 0x31, 0x25,
	0x2C, 0x06, 0x35, 0x04, 0x00, 0x2F, 0x31, 0x43, 0x51, 0x3B, 0x2E, 0x06,
	0x54, 0x55, 0x23, 0x18, 0x7A, 0x16, 0x2C, 0x57, 0x38, 0x7B, 0x18, 0x4E,
	0x3F, 0x2D, 0x21, 0x1D, 0x0C, 0x2F, 0x19, 0x14, 0x19, 0x22, 0x1B, 0x44,
	0x11, 0x0A, 0x32, 0x39, 0x2F, 0x31, 0x26, 0x1B, 0x02, 0x25, 0x0C, 0x2E,
	0x0E, 0x3A, 0x52, 0x09, 0x26, 0x0B, 0x27, 0x0E, 0x21, 0x3F, 0x31, 0x01,
	0x2A, 0x13, 0x59, 0x07, 0x23, 0x07, 0x18, 0x03, 0x50, 0x3C, 0x1F, 0x76,
	0x05, 0x33, 0x26, 0x53, 0x6D, 0x1E, 0x0C, 0x3E, 0x20, 0x10, 0x5E, 0x13,
	0x59, 0x18, 0x37, 0x23, 0x50, 0x5C, 0x05, 0x2C, 0x54, 0x56, 0x28, 0x52,
	0x34, 0x43, 0x3B, 0x37, 0x02, 0x2A, 0x26, 0x00, 0x3F, 0x2F, 0x35, 0x16,
	0x26, 0x28, 0x18, 0x17, 0x3E, 0x50, 0x25, 0x32, 0x15, 0x0E, 0x14, 0x38,
	0x24, 0x13, 0x25, 0x14, 0x1D, 0x5B, 0x04, 0x20, 0x55, 0x1C, 0x28, 0x01,
	0x2E, 0x08, 0x0F, 0x40, 0x08, 0x25, 0x0C, 0x1B, 0x40, 0x03, 0x23, 0x58,
	0x09, 0x19, 0x74, 0x14, 0x2E, 0x3C, 0x58, 0x0E, 0x0A, 0x09, 0x3D, 0x2E,
	0x38, 0x55, 0x56, 0x21, 0x03, 0x2C, 0x04, 0x0B, 0x2A, 0x22, 0x2D, 0x5F,
	0x19, 0x05, 0x27, 0x7B, 0x43, 0x25, 0x29, 0x13, 0x28, 0x2B, 0x28, 0x1F,
	0x07, 0x7A, 0x01, 0x15, 0x25, 0x58, 0x38, 0x43, 0x51, 0x01, 0x23, 0x73,
	0x0B, 0x31, 0x18, 0x09, 0x0F, 0x08, 0x3B, 0x5D, 0x02, 0x0D, 0x54, 0x3B,
	0x14, 0x08, 0x28, 0x5A, 0x32, 0x57, 0x22, 0x18, 0x5A, 0x4A, 0x57, 0x25,
	0x07, 0x2F, 0x2E, 0x2A, 0x5F, 0x70, 0x26, 0x24, 0x1F, 0x11, 0x6D, 0x08,
	0x0F, 0x41, 0x31, 0x12, 0x15, 0x57, 0x23, 0x52, 0x74, 0x3B, 0x07, 0x22,
	0x04, 0x3B, 0x24, 0x58, 0x2D, 0x38, 0x72, 0x47, 0x29, 0x0F, 0x1F, 0x23,
	0x58, 0x0C, 0x1E, 0x03, 0x0F, 0x21, 0x12, 0x36, 0x38, 0x13, 0x47, 0x52,
	0x3B, 0x1A, 0x03, 0x5F, 0x24, 0x01, 0x1A, 0x0E, 0x00, 0x39, 0x0B, 0x06,
	0x06, 0x3E, 0x30, 0x36, 0x52, 0x23, 0x22, 0x08, 0x19, 0x1D, 0x0F, 0x15,
	0x2C, 0x5A, 0x00, 0x0E, 0x19, 0x37, 0x28, 0x1E, 0x0A, 0x3E, 0x04, 0x02,
	0x22, 0x70, 0x3F, 0x0E, 0x20, 0x5A, 0x32, 0x5F, 0x06, 0x34, 0x01, 0x70,
	0x08, 0x0E, 0x18, 0x02, 0x2F, 0x1E, 0x0D, 0x34, 0x1C, 0x00, 0x23, 0x31,
	0x5B, 0x07, 0x30, 0x21, 0x38, 0x18, 0x3D, 0x14, 0x36, 0x06, 0x21, 0x5C,
	0x10, 0x54, 0x33, 0x1F, 0x1B, 0x32, 0x22, 0x26, 0x28, 0x01, 0x12, 0x00,
	0x23, 0x3A, 0x20, 0x35, 0x18, 0x35, 0x20, 0x2D, 0x75, 0x5B, 0x37, 0x34,
	0x44, 0x20, 0x5D, 0x36, 0x25, 0x44, 0x28, 0x04, 0x17, 0x5B, 0x24, 0x12,
	0x00, 0x4A, 0x1C, 0x2D, 0x75, 0x2F, 0x25, 0x21, 0x59, 0x16, 0x38, 0x34,
	0x01, 0x20, 0x7B, 0x59, 0x2C, 0x07, 0x00, 0x20, 0x3C, 0x33, 0x5E, 0x33,
	0x01, 0x38, 0x0A, 0x24, 0x02, 0x23, 0x1A, 0x58, 0x1A, 0x08, 0x28, 0x07,
	0x54, 0x5A, 0x39, 0x00, 0x59, 0x54, 0x25, 0x0D, 0x14, 0x3C, 0x10, 0x1A,
	0x21, 0x01, 0x06, 0x2E, 0x20, 0x33, 0x16, 0x39, 0x25, 0x1B, 0x2D, 0x0E,
	0x5B, 0x54, 0x2D, 0x09, 0x33, 0x0A, 0x23, 0x3A, 0x5D, 0x14, 0x38, 0x05,
	0x05, 0x12, 0x24, 0x38, 0x0C, 0x0F, 0x01, 0x35, 0x0D, 0x23, 0x1B, 0x5D,
	0x00, 0x16, 0x35, 0x0C, 0x3C, 0x0E, 0x58, 0x4E, 0x0D, 0x3B, 0x0B, 0x1A,
	0x18, 0x0F, 0x3F, 0x0E, 0x1A, 0x55, 0x3D, 0x59, 0x0F, 0x43, 0x36, 0x5D,
	0x58, 0x20, 0x55, 0x56, 0x45, 0x25, 0x10, 0x47, 0x0E, 0x1C, 0x52, 0x24,
	0x00, 0x09, 0x1C, 0x1D, 0x1A, 0x1B, 0x0C, 0x1E, 0x1B, 0x24, 0x3F, 0x0F,
	0x0A, 0x00, 0x7A, 0x3C, 0x37, 0x16, 0x07, 0x24, 0x1C, 0x2C, 0x3B, 0x19,
	0x03, 0x43, 0x0B, 0x39, 0x3D, 0x77, 0x39, 0x58, 0x45, 0x3F, 0x0E, 0x3B,
	0x4A, 0x0F, 0x05, 0x06, 0x1E, 0x59, 0x3F, 0x2F, 0x25, 0x19, 0x2D, 0x0C,
	0x3D, 0x20, 0x02, 0x39, 0x36, 0x22, 0x1B, 0x1D, 0x51, 0x57, 0x1F, 0x34,
	0x59, 0x04, 0x22, 0x19, 0x30, 0x18, 0x20, 0x56, 0x39, 0x71, 0x5A, 0x1B,
	0x39, 0x3B, 0x17, 0x3D, 0x2E, 0x03, 0x2F, 0x08, 0x3C, 0x51, 0x34, 0x0D,
	0x2B, 0x19, 0x12, 0x36, 0x53, 0x00, 0x3A, 0x30, 0x23, 0x32, 0x2D, 0x3F,
	0x36, 0x28, 0x0D, 0x1A, 0x20, 0x16, 0x2D, 0x22, 0x09, 0x43, 0x56, 0x0F,
	0x59, 0x3A, 0x43, 0x0D, 0x41, 0x0A, 0x10, 0x29, 0x17, 0x37, 0x3F, 0x2B,
	0x0E, 0x34, 0x24, 0x27, 0x18, 0x3B, 0x50, 0x5A, 0x19, 0x3B, 0x5A, 0x02,
	0x1A, 0x06, 0x29, 0x0A, 0x0F, 0x19, 0x22, 0x04, 0x5B, 0x22, 0x3E, 0x00,
	0x06, 0x3B, 0x11, 0x01, 0x1E, 0x21, 0x5E, 0x57, 0x2D, 0x12, 0x32, 0x3D,
	0x27, 0x34, 0x12, 0x28, 0x1B, 0x50, 0x2A, 0x5A, 0x2D, 0x2E, 0x23, 0x2C,
	0x18, 0x38, 0x5D, 0x0A, 0x07, 0x12, 0x31, 0x1E, 0x0E, 0x24, 0x1A, 0x1B,
	0x5C, 0x37, 0x41, 0x24, 0x3A, 0x0B, 0x2B, 0x2C, 0x1E, 0x16, 0x2A, 0x2F,
	0x5D, 0x23, 0x25, 0x20, 0x50, 0x02, 0x2E, 0x11, 0x5D, 0x23, 0x2B, 0x59,
	0x36, 0x2E, 0x0D, 0x0A, 0x44, 0x33, 0x3F, 0x29, 0x2B, 0x18, 0x24, 0x27,
	0x20, 0x0B, 0x24, 0x2A, 0x5D, 0x33, 0x3F, 0x09, 0x06, 0x55, 0x27, 0x24,
	0x28, 0x05, 0x00, 0x0C, 0x21, 0x09, 0x27, 0x1F, 0x19, 0x18, 0x5F, 0x21,
	0x2E, 0x26, 0x5D, 0x2E, 0x12, 0x5E, 0x34, 0x28, 0x5F, 0x09, 0x5D, 0x4A,
	0x19, 0x3A, 0x03, 0x0A, 0x58, 0x06, 0x1F, 0x1A, 0x0B, 0x31, 0x27, 0x44,
	0x0A, 0x06, 0x12, 0x2F, 0x06, 0x2D, 0x34, 0x31, 0x09, 0x5C, 0x10, 0x1B,
	0x32, 0x3C, 0x40, 0x12, 0x3D, 0x12, 0x07, 0x52, 0x0B, 0x21, 0x22, 0x41,
	0x39, 0x10, 0x0E, 0x30, 0x29, 0x5D, 0x06, 0x47, 0x0A, 0x18, 0x5C, 0x33,
	0x3C, 0x58, 0x07, 0x2D, 0x3A, 0x34, 0x29, 0x25, 0x32, 0x27, 0x43, 0x33,
	0x34, 0x2D, 0x24, 0x1B, 0x02, 0x2A, 0x20, 0x35, 0x0B, 0x2C, 0x16, 0x2C,
	0x2A, 0x28, 0x38, 0x38, 0x23, 0x34, 0x2D, 0x24, 0x0A, 0x44, 0x2F, 0x5D,
	0x2F, 0x2D, 0x2F, 0x03, 0x0D, 0x2D, 0x2A, 0x02, 0x7B, 0x47, 0x09, 0x08,
	0x2A, 0x2C, 0x1E, 0x39, 0x3F, 0x0A, 0x2B, 0x27, 0x34, 0x17, 0x02, 0x0F,
	0x54, 0x2A, 0x24, 0x08, 0x07, 0x02, 0x33, 0x0A, 0x2C, 0x16, 0x3E, 0x2E,
	0x2A, 0x2A, 0x12, 0x2E, 0x33, 0x58, 0x0A, 0x70, 0x1B, 0x31, 0x3E, 0x0A,
	0x07, 0x59, 0x20, 0x5C, 0x05, 0x16, 0x54, 0x55, 0x07, 0x07, 0x10, 0x58,
	0x14, 0x29, 0x2E, 0x12, 0x39, 0x23, 0x2B, 0x19, 0x0C, 0x36, 0x08, 0x27,
	0x5E, 0x2E, 0x3E, 0x0F, 0x38, 0x04, 0x04, 0x54, 0x29, 0x2D, 0x0A, 0x3B,
	0x24, 0x50, 0x0D, 0x21, 0x2A, 0x01, 0x0A, 0x09, 0x03, 0x0C, 0x20, 0x0A,
	0x27, 0x2A, 0x11, 0x0B, 0x54, 0x5C, 0x2F, 0x0A, 0x0D, 0x07, 0x5D, 0x20,
	0x12, 0x01, 0x12, 0x14, 0x1D, 0x0D, 0x47, 0x22, 0x3B, 0x02, 0x0F, 0x3C,
	0x56, 0x21, 0x1C, 0x03, 0x3E, 0x02, 0x05, 0x5E, 0x37, 0x01, 0x2F, 0x0F,
	0x08, 0x30, 0x35, 0x31, 0x23, 0x01, 0x08, 0x22, 0x39, 0x1C, 0x0F, 0x74,
	0x2F, 0x09, 0x1D, 0x27, 0x29, 0x04, 0x56, 0x56, 0x2F, 0x7B, 0x1D, 0x29,
	0x3E, 0x01, 0x31, 0x3F, 0x4A, 0x5F, 0x00, 0x06, 0x2B, 0x50, 0x38, 0x3B,
	0x0F, 0x3E, 0x05, 0x1C, 0x26, 0x0B, 0x2D, 0x55, 0x05, 0x3A, 0x2B, 0x38,
	0x4E, 0x36, 0x5F, 0x0B, 0x27, 0x02, 0x0B, 0x22, 0x2A, 0x5B, 0x27, 0x34,
	0x5D, 0x0A, 0x04, 0x23, 0x28, 0x52, 0x04, 0x35, 0x55, 0x56, 0x52, 0x7A,
	0x28, 0x58, 0x39, 0x5B, 0x0B, 0x2A, 0x22, 0x0C, 0x1A, 0x11, 0x55, 0x36,
	0x3F, 0x2D, 0x0B, 0x2B, 0x06, 0x3D, 0x59, 0x3B, 0x19, 0x11, 0x36, 0x3D,
	0x0C, 0x25, 0x57, 0x59, 0x53, 0x13, 0x14, 0x36, 0x01, 0x09, 0x0E, 0x23,
	0x08, 0x28, 0x5B, 0x10, 0x1C, 0x59, 0x01, 0x5B, 0x2B, 0x36, 0x20, 0x41,
	0x04, 0x74, 0x2E, 0x23, 0x22, 0x20, 0x2A, 0x2B, 0x0F, 0x58, 0x23, 0x0E,
	0x02, 0x1B, 0x36, 0x0C, 0x0B, 0x1B, 0x03, 0x38, 0x18, 0x2B, 0x2E, 0x59,
	0x1C, 0x24, 0x34, 0x43, 0x12, 0x26, 0x52, 0x26, 0x5D, 0x33, 0x3F, 0x59,
	0x37, 0x36, 0x50, 0x0A, 0x58, 0x14, 0x58, 0x53, 0x3C, 0x06, 0x74, 0x5B,
	0x30, 0x3A, 0x2E, 0x09, 0x0E, 0x0C, 0x26, 0x09, 0x28, 0x39, 0x0E, 0x29,
	0x0F, 0x03, 0x2E, 0x2B, 0x3F, 0x18, 0x7A, 0x03, 0x52, 0x1F, 0x19, 0x14,
	0x47, 0x20, 0x03, 0x29, 0x0A, 0x2D, 0x34, 0x5A, 0x44, 0x23, 0x18, 0x1B,
	0x0D, 0x33, 0x76, 0x24, 0x31, 0x14, 0x5E, 0x7B, 0x3F, 0x32, 0x2D, 0x0C,
	0x0E, 0x1B, 0x0F, 0x2F, 0x25, 0x01, 0x1A, 0x05, 0x27, 0x3C, 0x3B, 0x38,
	0x53, 0x0D, 0x33, 0x72, 0x3D, 0x08, 0x1B, 0x3A, 0x76, 0x2B, 0x19, 0x27,
	0x28, 0x0E, 0x28, 0x20, 0x2A, 0x59, 0x09, 0x2E, 0x2F, 0x3F, 0x06, 0x00,
	0x03, 0x37, 0x04, 0x0C, 0x37, 0x03, 0x35, 0x2F, 0x3F, 0x6D, 0x2D, 0x54,
	0x58, 0x2C, 0x21, 0x20, 0x2C, 0x1D, 0x22, 0x70, 0x04, 0x19, 0x2F, 0x3E,
	0x15, 0x01, 0x29, 0x21, 0x01, 0x73, 0x36, 0x03, 0x3D, 0x0C, 0x20, 0x01,
	0x4E, 0x2F, 0x3D, 0x29, 0x43, 0x2F, 0x39, 0x5E, 0x74, 0x2F, 0x26, 0x37,
	0x33, 0x29, 0x20, 0x59, 0x5C, 0x04, 0x16, 0x58, 0x55, 0x38, 0x02, 0x2B,
	0x5A, 0x18, 0x05, 0x3A, 0x13, 0x1E, 0x57, 0x03, 0x2E, 0x0A, 0x06, 0x2D,
	0x5A, 0x19, 0x6D, 0x27, 0x55, 0x1F, 0x18, 0x08, 0x54, 0x35, 0x0D, 0x00,
	0x3A, 0x28, 0x59, 0x0D, 0x02, 0x73, 0x47, 0x39, 0x2B, 0x29, 0x2B, 0x26,
	0x23, 0x0C, 0x5D, 0x14, 0x29, 0x31, 0x06, 0x0F, 0x0E, 0x20, 0x20, 0x45,
	0x22, 0x20, 0x2D, 0x56, 0x28, 0x19, 0x25, 0x59, 0x58, 0x18, 0x00, 0x24,
	0x27, 0x2C, 0x3F, 0x1B, 0x20, 0x2F, 0x2E, 0x2B, 0x2F, 0x21, 0x1E, 0x2C,
	0x3F, 0x04, 0x07, 0x0E, 0x11, 0x5B, 0x20, 0x0A, 0x18, 0x2A, 0x1F, 0x01,
	0x05, 0x38, 0x30, 0x0D, 0x0A, 0x0B, 0x59, 0x35, 0x0D, 0x3F, 0x73, 0x24,
	0x4E, 0x05, 0x0C, 0x0D, 0x0D, 0x14, 0x25, 0x31, 0x0A, 0x47, 0x52, 0x1A,
	0x2A, 0x2C, 0x3D, 0x50, 0x37, 0x2E, 0x05, 0x39, 0x2B, 0x3C, 0x27, 0x23,
	0x3B, 0x27, 0x02, 0x2F, 0x0C, 0x29, 0x03, 0x04, 0x18, 0x25, 0x2E, 0x2C,
	0x27, 0x3A, 0x27, 0x38, 0x39, 0x5B, 0x21, 0x7A, 0x2F, 0x27, 0x06, 0x5D,
	0x0A, 0x05, 0x51, 0x56, 0x2F, 0x00, 0x2E, 0x26, 0x01, 0x59, 0x09, 0x01,
	0x29, 0x09, 0x3C, 0x25, 0x1D, 0x27, 0x05, 0x09, 0x23, 0x35, 0x38, 0x01,
	0x28, 0x11, 0x24, 0x30, 0x23, 0x28, 0x13, 0x59, 0x57, 0x2C, 0x20, 0x2C,
	0x5B, 0x52, 0x2F, 0x27, 0x13, 0x3F, 0x0F, 0x08, 0x01, 0x27, 0x5B, 0x2E,
	0x5E, 0x40, 0x28, 0x1B, 0x33, 0x5F, 0x40, 0x23, 0x19, 0x31, 0x27, 0x29,
	0x0C, 0x27, 0x2D, 0x25, 0x27, 0x7A, 0x19, 0x50, 0x07, 0x28, 0x34, 0x01,
	0x26, 0x0D, 0x06, 0x05, 0x1B, 0x2A, 0x5F, 0x22, 0x25, 0x02, 0x05, 0x41,
	0x25, 0x71, 0x2B, 0x0A, 0x1E, 0x2F, 0x35, 0x0F, 0x05, 0x3D, 0x1D, 0x05,
	0x22, 0x2C, 0x05, 0x09, 0x12, 0x3A, 0x58, 0x0D, 0x40, 0x10, 0x0B, 0x16,
	0x37, 0x03, 0x04, 0x09, 0x53, 0x28, 0x2A, 0x70, 0x3F, 0x2B, 0x45, 0x03,
	0x11, 0x1F, 0x10, 0x1D, 0x19, 0x06, 0x3F, 0x52, 0x18, 0x2A, 0x26, 0x55,
	0x59, 0x0D, 0x02, 0x0C, 0x0E, 0x12, 0x39, 0x3D, 0x01, 0x1F, 0x25, 0x02,
	0x5C, 0x13, 0x2B, 0x27, 0x41, 0x23, 0x18, 0x39, 0x0C, 0x18, 0x59, 0x06,
	0x26, 0x26, 0x56, 0x01, 0x3A, 0x2D, 0x55, 0x2D, 0x00, 0x13, 0x1F, 0x0A,
	0x0D, 0x0E, 0x0D, 0x3F, 0x16, 0x5C, 0x01, 0x30, 0x3E, 0x16, 0x0B, 0x0F,
	0x1B, 0x3E, 0x11, 0x56, 0x03, 0x2C, 0x59, 0x23, 0x3A, 0x0D, 0x05, 0x58,
	0x59, 0x1C, 0x1F, 0x2A, 0x1A, 0x15, 0x14, 0x06, 0x08, 0x27, 0x29, 0x09,
	0x2E, 0x2C, 0x36, 0x22, 0x18, 0x1B, 0x15, 0x0E, 0x1B, 0x56, 0x28, 0x25,
	0x43, 0x54, 0x2C, 0x31, 0x7A, 0x1B, 0x54, 0x25, 0x1E, 0x00, 0x43, 0x51,
	0x3B, 0x27, 0x09, 0x58, 0x2C, 0x3F, 0x58, 0x2F, 0x3E, 0x59, 0x00, 0x2A,
	0x3A, 0x21, 0x0A, 0x19, 0x5E, 0x71, 0x20, 0x55, 0x0C, 0x01, 0x25, 0x28,
	0x31, 0x20, 0x5B, 0x0A, 0x1A, 0x52, 0x5D, 0x1C, 0x05, 0x58, 0x39, 0x08,
	0x1A, 0x0E, 0x0F, 0x52, 0x58, 0x0A, 0x04, 0x08, 0x11, 0x20, 0x0A, 0x0F,
	0x23, 0x0E, 0x28, 0x38, 0x72, 0x0B, 0x16, 0x3A, 0x27, 0x27, 0x16, 0x2C,
	0x5B, 0x38, 0x03, 0x1D, 0x56, 0x3F, 0x27, 0x0D, 0x1F, 0x34, 0x2D, 0x3D,
	0x26, 0x3D, 0x0D, 0x20, 0x3C, 0x36, 0x55, 0x19, 0x29, 0x21, 0x00, 0x3E,
	0x30, 0x3F, 0x2F, 0x3A, 0x0D, 0x34, 0x3A, 0x23, 0x18, 0x38, 0x35, 0x25,
	0x0A, 0x07, 0x22, 0x31, 0x5A, 0x2D, 0x09, 0x22, 0x05, 0x07, 0x24, 0x0B,
	0x5E, 0x2A, 0x5A, 0x3A, 0x21, 0x5E, 0x0F, 0x36, 0x06, 0x26, 0x3F, 0x27,
	0x06, 0x19, 0x26, 0x19, 0x14, 0x3B, 0x25, 0x74, 0x5D, 0x06, 0x26, 0x0F,
	0x10, 0x55, 0x11, 0x5B, 0x12, 0x0C, 0x1F, 0x09, 0x3D, 0x2E, 0x32, 0x3A,
	0x34, 0x1D, 0x3D, 0x25, 0x34, 0x02, 0x2A, 0x02, 0x03, 0x07, 0x2B, 0x09,
	0x59, 0x15, 0x5B, 0x15, 0x0A, 0x31, 0x16, 0x55, 0x12, 0x00, 0x1B, 0x37,
	0x5B, 0x36, 0x24, 0x1B, 0x74, 0x1F, 0x22, 0x1E, 0x59, 0x26, 0x03, 0x14,
	0x26, 0x2A, 0x0D, 0x5E, 0x00, 0x04, 0x0F, 0x72, 0x14, 0x07, 0x14, 0x04,
	0x33, 0x34, 0x30, 0x3B, 0x0C, 0x13, 0x35, 0x37, 0x17, 0x27, 0x09, 0x58,
	0x00, 0x03, 0x26, 0x34, 0x36, 0x00, 0x0C, 0x53, 0x3A, 0x25, 0x59, 0x21,
	0x3A, 0x30, 0x08, 0x20, 0x1B, 0x11, 0x34, 0x09, 0x28, 0x17, 0x3D, 0x25,
	0x58, 0x0F, 0x28, 0x5B, 0x2E, 0x0D, 0x23, 0x1F, 0x3A, 0x75, 0x59, 0x29,
	0x2A, 0x00, 0x0C, 0x3B, 0x2E, 0x56, 0x5B, 0x29, 0x0F, 0x02, 0x3A, 0x1B,
	0x15, 0x5E, 0x4E, 0x2B, 0x3A, 0x13, 0x5F, 0x24, 0x0D, 0x31, 0x33, 0x3B,
	0x52, 0x2B, 0x24, 0x08, 0x0E, 0x34, 0x27, 0x11, 0x2D, 0x0B, 0x29, 0x2A,
	0x3E, 0x3A, 0x2E, 0x35, 0x0C, 0x25, 0x15, 0x3B, 0x0F, 0x5C, 0x3F, 0x10,
	0x3D, 0x32, 0x3D, 0x01, 0x1B, 0x23, 0x54, 0x22, 0x0D, 0x10, 0x28, 0x3B,
	0x0C, 0x3C, 0x2C, 0x3B, 0x36, 0x0F, 0x1F, 0x20, 0x54, 0x39, 0x3B, 0x1F,
	0x04, 0x25, 0x12, 0x59, 0x1C, 0x73, 0x26, 0x39, 0x17, 0x2F, 0x14, 0x5A,
	0x08, 0x16, 0x09, 0x7A, 0x28, 0x10, 0x23, 0x5C, 0x3A, 0x25, 0x50, 0x0C,
	0x53, 0x05, 0x1A, 0x0A, 0x5D, 0x18, 0x28, 0x54, 0x17, 0x36, 0x5D, 0x2A,
	0x08, 0x06, 0x29, 0x1E, 0x7B, 0x01, 0x52, 0x3A, 0x1F, 0x2A, 0x16, 0x39,
	0x3D, 0x3F, 0x74, 0x04, 0x25, 0x2D, 0x59, 0x01, 0x2B, 0x2D, 0x1E, 0x2A,
	0x3A, 0x08, 0x18, 0x0B, 0x2A, 0x00, 0x3A, 0x1B, 0x5C, 0x02, 0x2D, 0x0F,
	0x0A, 0x18, 0x09, 0x06, 0x2F, 0x20, 0x24, 0x3E, 0x70, 0x3B, 0x3B, 0x05,
	0x28, 0x3A, 0x04, 0x2B, 0x3B, 0x2D, 0x38, 0x5B, 0x37, 0x03, 0x0E, 0x28,
	0x3D, 0x2F, 0x37, 0x1A, 0x2D, 0x3B, 0x3B, 0x01, 0x1D, 0x27, 0x1B, 0x0B,
	0x16, 0x39, 0x0F, 0x2E, 0x2B, 0x1A, 0x21, 0x75, 0x39, 0x55, 0x45, 0x5A,
	0x0E, 0x5E, 0x29, 0x1D, 0x13, 0x0E, 0x19, 0x50, 0x02, 0x5B, 0x0C, 0x02,
	0x07, 0x29, 0x52, 0x09, 0x3A, 0x0D, 0x5A, 0x5C, 0x74, 0x3B, 0x50, 0x21,
	0x13, 0x13, 0x04, 0x02, 0x5C, 0x07, 0x09, 0x09, 0x06, 0x3C, 0x32, 0x3B,
	0x58, 0x12, 0x34, 0x5A, 0x3A, 0x05, 0x0A, 0x5A, 0x5D, 0x0F, 0x1F, 0x33,
	0x03, 0x1E, 0x72, 0x58, 0x09, 0x2A, 0x5E, 0x08, 0x3B, 0x34, 0x5F, 0x29,
	0x0C, 0x21, 0x27, 0x39, 0x27, 0x75, 0x55, 0x04, 0x37, 0x22, 0x09, 0x0F,
	0x2B, 0x04, 0x03, 0x76, 0x15, 0x20, 0x28, 0x2D, 0x33, 0x5F, 0x58, 0x14,
	0x19, 0x2A, 0x5E, 0x27, 0x18, 0x59, 0x09, 0x0F, 0x35, 0x2F, 0x3B, 0x03,
	0x02, 0x12, 0x26, 0x32, 0x2B, 0x15, 0x2B, 0x07, 0x3D, 0x27, 0x00, 0x06,
	0x5F, 0x1E, 0x1A, 0x1A, 0x51, 0x1B, 0x44, 0x0A, 0x38, 0x04, 0x17, 0x07,
	0x72, 0x2A, 0x30, 0x04, 0x3C, 0x01, 0x1F, 0x2E, 0x1C, 0x23, 0x0D, 0x5F,
	0x15, 0x0A, 0x5B, 0x2E, 0x3D, 0x56, 0x38, 0x1D, 0x2F, 0x03, 0x33, 0x0F,
	0x3A, 0x10, 0x25, 0x0B, 0x0D, 0x08, 0x2E, 0x22, 0x54, 0x5F, 0x22, 0x21,
	0x0F, 0x27, 0x0A, 0x21, 0x69, 0x1B, 0x0E, 0x1F, 0x11, 0x70, 0x5E, 0x27,
	0x39, 0x3D, 0x2B, 0x1B, 0x4E, 0x04, 0x27, 0x07, 0x28, 0x51, 0x36, 0x5B,
	0x1B, 0x3A, 0x06, 0x3E, 0x3F, 0x05, 0x3A, 0x10, 0x1F, 0x3B, 0x18, 0x1E,
	0x05, 0x20, 0x26, 0x01, 0x2F, 0x10, 0x3C, 0x5E, 0x2D, 0x2D, 0x2D, 0x5B,
	0x23, 0x2D, 0x1F, 0x2E, 0x0C, 0x5E, 0x00, 0x58, 0x23, 0x25, 0x32, 0x35,
	0x05, 0x34, 0x18, 0x03, 0x24, 0x28, 0x53, 0x28, 0x3E, 0x10, 0x05, 0x2E,
	0x57, 0x0E, 0x01, 0x03, 0x31, 0x27, 0x02, 0x33, 0x0B, 0x10, 0x21, 0x12,
	0x28, 0x5D, 0x19, 0x26, 0x3D, 0x14, 0x5D, 0x55, 0x2F, 0x0C, 0x73, 0x3E,
	0x37, 0x05, 0x31, 0x32, 0x5B, 0x1B, 0x5D, 0x05, 0x34, 0x2B, 0x13, 0x2C,
	0x1C, 0x00, 0x3F, 0x29, 0x5F, 0x3F, 0x06, 0x07, 0x2E, 0x18, 0x5A, 0x1A,
	0x07, 0x58, 0x1F, 0x2A, 0x09, 0x1F, 0x2E, 0x59, 0x20, 0x23, 0x3D, 0x18,
	0x1C, 0x25, 0x2B, 0x0D, 0x10, 0x01, 0x40, 0x0A, 0x5E, 0x17, 0x02, 0x0F,
	0x08, 0x24, 0x10, 0x3D, 0x13, 0x08, 0x3A, 0x1B, 0x56, 0x2F, 0x01, 0x27,
	0x02, 0x1B, 0x18, 0x18, 0x0E, 0x4A, 0x56, 0x2E, 0x21, 0x09, 0x34, 0x02,
	0x1A, 0x05, 0x3D, 0x11, 0x20, 0x5A, 0x35, 0x1C, 0x36, 0x37, 0x24, 0x11,
	0x18, 0x4A, 0x0A, 0x24, 0x21, 0x3F, 0x39, 0x0B, 0x02, 0x26, 0x24, 0x16,
	0x5C, 0x01, 0x6D, 0x47, 0x59, 0x37, 0x53, 0x2B, 0x36, 0x39, 0x01, 0x12,
	0x27, 0x1A, 0x2B, 0x3C, 0x33, 0x15, 0x06, 0x55, 0x41, 0x00, 0x1B, 0x0E,
	0x14, 0x18, 0x09, 0x32, 0x14, 0x0B, 0x56, 0x23, 0x77, 0x06, 0x0F, 0x2B,
	0x39, 0x20, 0x1A, 0x0C, 0x07, 0x3A, 0x37, 0x43, 0x33, 0x0F, 0x08, 0x69,
	0x20, 0x4E, 0x02, 0x1C, 0x6D, 0x5B, 0x58, 0x5E, 0x24, 0x6D, 0x16, 0x11,
	0x17, 0x5D, 0x38, 0x5E, 0x51, 0x0B, 0x3C, 0x00, 0x03, 0x54, 0x38, 0x28,
	0x74, 0x27, 0x2C, 0x0B, 0x00, 0x00, 0x23, 0x15, 0x03, 0x26, 0x0B, 0x26,
	0x0C, 0x20, 0x5B, 0x76, 0x0B, 0x10, 0x01, 0x39, 0x2D, 0x04, 0x19, 0x28,
	0x05, 0x72, 0x2F, 0x31, 0x2F, 0x52, 0x14, 0x22, 0x08, 0x1A, 0x23, 0x37,
	0x2F, 0x0E, 0x0F, 0x25, 0x10, 0x0F, 0x2B, 0x1B, 0x2E, 0x04, 0x39, 0x53,
	0x5B, 0x18, 0x2E, 0x02, 0x59, 0x3D, 0x08, 0x37, 0x0E, 0x58, 0x2C, 0x59,
	0x31, 0x07, 0x23, 0x0D, 0x5C, 0x07, 0x20, 0x07, 0x3E, 0x07, 0x7B, 0x2D,
	0x0A, 0x06, 0x40, 0x28, 0x08, 0x18, 0x2F, 0x26, 0x21, 0x39, 0x35, 0x19,
	0x5C, 0x7A, 0x5C, 0x09, 0x19, 0x2E, 0x27, 0x08, 0x38, 0x02, 0x31, 0x2A,
	0x2B, 0x31, 0x59, 0x53, 0x0B, 0x0B, 0x33, 0x41, 0x1B, 0x29, 0x3A, 0x02,
	0x45, 0x0A, 0x0A, 0x15, 0x35, 0x3F, 0x5D, 0x72, 0x08, 0x30, 0x5B, 0x23,
	0x2C, 0x24, 0x2D, 0x04, 0x3F, 0x01, 0x34, 0x25, 0x2A, 0x00, 0x0E, 0x19,
	0x27, 0x19, 0x33, 0x15, 0x06, 0x51, 0x2D, 0x08, 0x37, 0x35, 0x36, 0x57,
	0x58, 0x34, 0x5C, 0x08, 0x07, 0x2C, 0x23, 0x14, 0x57, 0x04, 0x22, 0x17,
	0x0D, 0x23, 0x18, 0x3F, 0x01, 0x1C, 0x30, 0x26, 0x11, 0x6D, 0x0B, 0x26,
	0x09, 0x0F, 0x03, 0x3F, 0x07, 0x27, 0x3E, 0x76, 0x20, 0x08, 0x08, 0x5E,
	0x01, 0x1C, 0x2F, 0x37, 0x11, 0x24, 0x15, 0x30, 0x04, 0x0C, 0x10, 0x3F,
	0x02, 0x01, 0x2D, 0x11, 0x5E, 0x14, 0x1D, 0x19, 0x00, 0x25, 0x0A, 0x00,
	0x2C, 0x1A, 0x5E, 0x27, 0x3C, 0x1D, 0x25, 0x14, 0x4A, 0x3F, 0x1B, 0x0C,
	0x06, 0x2E, 0x3F, 0x2F, 0x10, 0x1C, 0x28, 0x2D, 0x21, 0x04, 0x5E, 0x4A,
	0x19, 0x03, 0x10, 0x58, 0x35, 0x3E, 0x3E, 0x14, 0x1C, 0x12, 0x24, 0x3B,
	0x2F, 0x1D, 0x59, 0x19, 0x01, 0x18, 0x2B, 0x59, 0x19, 0x2E, 0x28, 0x3F,
	0x06, 0x0B, 0x3A, 0x75, 0x34, 0x53, 0x2B, 0x5D, 0x12, 0x2D, 0x56, 0x17,
	0x2D, 0x27, 0x20, 0x52, 0x2C, 0x1D, 0x31, 0x27, 0x23, 0x14, 0x24, 0x11,
	0x0B, 0x55, 0x19, 0x00, 0x03, 0x5C, 0x08, 0x21, 0x40, 0x35, 0x03, 0x1B,
	0x5A, 0x2F, 0x0A, 0x38, 0x37, 0x5B, 0x0C, 0x08, 0x3C, 0x51, 0x20, 0x53,
	0x2A, 0x39, 0x2C, 0x37, 0x12, 0x17, 0x36, 0x26, 0x27, 0x0C, 0x0E, 0x26,
	0x34, 0x38, 0x40, 0x2A, 0x2F, 0x28, 0x57, 0x06, 0x1A, 0x5A, 0x24, 0x34,
	0x0D, 0x30, 0x26, 0x59, 0x06, 0x3D, 0x2F, 0x21, 0x54, 0x2C, 0x21, 0x05,
	0x21, 0x09, 0x3C, 0x22, 0x0D, 0x02, 0x53, 0x28, 0x3A, 0x69, 0x2A, 0x19,
	0x03, 0x20, 0x7B, 0x1B, 0x26, 0x3E, 0x13, 0x29, 0x47, 0x16, 0x1F, 0x11,
	0x05, 0x0F, 0x0C, 0x1E, 0x25, 0x01, 0x20, 0x2B, 0x2F, 0x39, 0x0E, 0x3A,
	0x37, 0x5B, 0x0C, 0x06, 0x06, 0x4A, 0x08, 0x5E, 0x01, 0x1F, 0x4A, 0x2A,
	0x05, 0x6D, 0x22, 0x58, 0x06, 0x0E, 0x21, 0x16, 0x0A, 0x1B, 0x52, 0x16,
	0x05, 0x36, 0x3F, 0x5F, 0x29, 0x24, 0x1B, 0x04, 0x20, 0x3A, 0x1B, 0x2E,
	0x04, 0x13, 0x24, 0x58, 0x22, 0x07, 0x40, 0x03, 0x02, 0x19, 0x29, 0x40,
	0x35, 0x04, 0x26, 0x23, 0x31, 0x01, 0x1F, 0x0B, 0x1B, 0x39, 0x00, 0x25,
	0x2E, 0x00, 0x12, 0x04, 0x2A, 0x59, 0x22, 0x01, 0x11, 0x2A, 0x4E, 0x06,
	0x38, 0x12, 0x0B, 0x3B, 0x5B, 0x38, 0x31, 0x0F, 0x19, 0x3B, 0x01, 0x69,
	0x1B, 0x24, 0x09, 0x1E, 0x03, 0x1C, 0x2A, 0x18, 0x0D, 0x0B, 0x39, 0x39,
	0x19, 0x0E, 0x12, 0x2A, 0x17, 0x1D, 0x20, 0x0E, 0x58, 0x02, 0x08, 0x02,
	0x09, 0x5B, 0x30, 0x19, 0x00, 0x2C, 0x1F, 0x38, 0x17, 0x3C, 0x25, 0x0B,
	0x4A, 0x0A, 0x13, 0x1A, 0x23, 0x23, 0x01, 0x0E, 0x3A, 0x43, 0x06, 0x25,
	0x13, 0x7A, 0x28, 0x31, 0x39, 0x2D, 0x6D, 0x04, 0x36, 0x2B, 0x32, 0x3B,
	0x05, 0x3B, 0x26, 0x00, 0x03, 0x1F, 0x0A, 0x0B, 0x33, 0x70, 0x29, 0x14,
	0x3E, 0x22, 0x75, 0x16, 0x27, 0x37, 0x5D, 0x06, 0x02, 0x51, 0x1A, 0x53,
	0x2A, 0x36, 0x02, 0x19, 0x2E, 0x2A, 0x21, 0x0B, 0x1B, 0x39, 0x10, 0x25,
	0x05, 0x18, 0x00, 0x09, 0x20, 0x55, 0x36, 0x23, 0x7A, 0x0E, 0x56, 0x2D,
	0x53, 0x24, 0x2E, 0x0B, 0x57, 0x39, 0x14, 0x0D, 0x26, 0x0D, 0x06, 0x2C,
	0x27, 0x34, 0x3C, 0x12, 0x05, 0x0F, 0x18, 0x41, 0x21, 0x7A, 0x26, 0x16,
	0x20, 0x39, 0x04, 0x25, 0x05, 0x41, 0x04, 0x09, 0x20, 0x59, 0x3E, 0x03,
	0x3B, 0x00, 0x05, 0x5A, 0x24, 0x1B, 0x59, 0x36, 0x18, 0x18, 0x0B, 0x26,
	0x53, 0x07, 0x52, 0x00, 0x2B, 0x2F, 0x23, 0x32, 0x25, 0x54, 0x31, 0x22,
	0x1F, 0x73, 0x5F, 0x15, 0x20, 0x27, 0x2D, 0x0F, 0x0A, 0x5E, 0x19, 0x13,
	0x1F, 0x00, 0x5B, 0x58, 0x12, 0x43, 0x25, 0x18, 0x1E, 0x33, 0x1B, 0x57,
	0x27, 0x12, 0x72, 0x5B, 0x1B, 0x1F, 0x22, 0x3A, 0x1C, 0x0F, 0x5D, 0x31,
	0x0E, 0x07, 0x52, 0x1E, 0x13, 0x0F, 0x1F, 0x0C, 0x23, 0x21, 0x09, 0x38,
	0x19, 0x3F, 0x04, 0x77, 0x55, 0x26, 0x04, 0x3B, 0x3A, 0x01, 0x2B, 0x38,
	0x28, 0x11, 0x14, 0x36, 0x08, 0x2C, 0x16, 0x5A, 0x37, 0x24, 0x26, 0x75,
	0x0F, 0x30, 0x28, 0x03, 0x29, 0x20, 0x0B, 0x17, 0x3C, 0x01, 0x0A, 0x05,
	0x02, 0x1F, 0x1B, 0x3A, 0x06, 0x04, 0x5F, 0x3B, 0x3F, 0x29, 0x1E, 0x3C,
	0x0A, 0x54, 0x0A, 0x29, 0x5B, 0x2D, 0x1F, 0x18, 0x04, 0x19, 0x28, 0x09,
	0x17, 0x1D, 0x2D, 0x2B, 0x3A, 0x32, 0x2D, 0x29, 0x24, 0x3C, 0x22, 0x3E,
	0x00, 0x06, 0x55, 0x59, 0x03, 0x5C, 0x21, 0x1A, 0x30, 0x58, 0x11, 0x74,
	0x3D, 0x16, 0x24, 0x1B, 0x3A, 0x03, 0x4A, 0x3C, 0x33, 0x2D, 0x2B, 0x35,
	0x5E, 0x24, 0x30, 0x26, 0x05, 0x28, 0x28, 0x05, 0x07, 0x36, 0x37, 0x24,
	0x0B, 0x26, 0x52, 0x00, 0x58, 0x17, 0x15, 0x0A, 0x2C, 0x1F, 0x04, 0x34,
	0x51, 0x26, 0x05, 0x70, 0x38, 0x2B, 0x39, 0x3C, 0x08, 0x0A, 0x23, 0x5E,
	0x29, 0x00, 0x3D, 0x03, 0x1C, 0x09, 0x0C, 0x47, 0x12, 0x1A, 0x38, 0x24,
	0x0D, 0x07, 0x00, 0x23, 0x7B, 0x3A, 0x2A, 0x18, 0x04, 0x75, 0x22, 0x15,
	0x20, 0x21, 0x2D, 0x3C, 0x58, 0x04, 0x32, 0x2F, 0x59, 0x04, 0x56, 0x38,
	0x14, 0x5D, 0x35, 0x3D, 0x22, 0x20, 0x06, 0x15, 0x0B, 0x0C, 0x72, 0x2B,
	0x23, 0x0C, 0x00, 0x0C, 0x07, 0x0E, 0x22, 0x5B, 0x76, 0x1D, 0x0D, 0x5B,
	0x03, 0x25, 0x59, 0x28, 0x1C, 0x31, 0x17, 0x0A, 0x50, 0x36, 0x53, 0x74,
	0x20, 0x50, 0x14, 0x18, 0x38, 0x5B, 0x30, 0x5D, 0x01, 0x29, 0x3B, 0x0B,
	0x58, 0x20, 0x2E, 0x20, 0x2C, 0x38, 0x59, 0x75, 0x28, 0x2C, 0x37, 0x3D,
	0x27, 0x3F, 0x12, 0x1B, 0x00, 0x27, 0x2D, 0x0C, 0x28, 0x2D, 0x75, 0x22,
	0x0A, 0x09, 0x40, 0x0F, 0x2D, 0x23, 0x3E, 0x1D, 0x76, 0x14, 0x0E, 0x58,
	0x0A, 0x0B, 0x26, 0x09, 0x38, 0x02, 0x34, 0x2D, 0x28, 0x5D, 0x0D, 0x2B,
	0x35, 0x15, 0x20, 0x2F, 0x1A, 0x18, 0x16, 0x29, 0x12, 0x08, 0x02, 0x17,
	0x5F, 0x32, 0x21, 0x05, 0x2F, 0x22, 0x0D, 0x30, 0x24, 0x12, 0x22, 0x26,
	0x75, 0x18, 0x2A, 0x37, 0x2E, 0x38, 0x22, 0x35, 0x2D, 0x0F, 0x0E, 0x25,
	0x57, 0x5C, 0x03, 0x72, 0x07, 0x0B, 0x0F, 0x07, 0x74, 0x1A, 0x4A, 0x3F,
	0x32, 0x30, 0x0E, 0x20, 0x25, 0x24, 0x24, 0x1E, 0x17, 0x56, 0x1D, 0x72,
	0x34, 0x54, 0x41, 0x40, 0x69, 0x5A, 0x1B, 0x45, 0x40, 0x74, 0x1E, 0x4A,
	0x39, 0x5D, 0x6D, 0x43, 0x15, 0x1B, 0x1A, 0x6D, 0x19, 0x16, 0x36, 0x59,
	0x2A, 0x3F, 0x1B, 0x57, 0x28, 0x6D, 0x3C, 0x2B, 0x0B, 0x33, 0x24, 0x23,
	0x08, 0x3C, 0x3E, 0x01, 0x1A, 0x37, 0x34, 0x5A, 0x31, 0x01, 0x56, 0x57,
	0x2D, 0x75, 0x5D, 0x38, 0x5A, 0x1E, 0x7B, 0x1B, 0x4E, 0x36, 0x0E, 0x7A,
	0x43, 0x0B, 0x1A, 0x31, 0x6D, 0x5C, 0x36, 0x22, 0x20, 0x29, 0x15, 0x14,
	0x08, 0x3A, 0x14, 0x20, 0x13, 0x02, 0x3A, 0x12, 0x14, 0x59, 0x5F, 0x40,
	0x20, 0x3E, 0x07, 0x1E, 0x0A, 0x75, 0x22, 0x18, 0x22, 0x3F, 0x13, 0x09,
	0x03, 0x58, 0x33, 0x10, 0x02, 0x06, 0x5D, 0x3A, 0x05, 0x06, 0x38, 0x38,
	0x5D, 0x32, 0x06, 0x18, 0x26, 0x1E, 0x72, 0x3A, 0x0F, 0x2B, 0x44, 0x10,
	0x23, 0x34, 0x03, 0x5E, 0x2E, 0x5D, 0x0D, 0x17, 0x04, 0x07, 0x39, 0x16,
	0x00, 0x1E, 0x24, 0x3C, 0x03, 0x5B, 0x33, 0x07, 0x5A, 0x05, 0x1D, 0x07,
	0x18, 0x01, 0x1B, 0x38, 0x0F, 0x25, 0x05, 0x15, 0x59, 0x12, 0x11, 0x59,
	0x2D, 0x0F, 0x44, 0x7B, 0x1C, 0x2D, 0x06, 0x5F, 0x2B, 0x18, 0x0A, 0x06,
	0x31, 0x29, 0x5C, 0x3B, 0x2C, 0x06, 0x10, 0x01, 0x2A, 0x36, 0x52, 0x75,
	0x47, 0x33, 0x2B, 0x5B, 0x2F, 0x43, 0x3B, 0x5C, 0x52, 0x03, 0x2A, 0x2B,
	0x1D, 0x00, 0x34, 0x26, 0x26, 0x2D, 0x32, 0x08, 0x06, 0x04, 0x14, 0x5F,
	0x77, 0x14, 0x52, 0x01, 0x5F, 0x7A, 0x03, 0x4E, 0x38, 0x21, 0x09, 0x16,
	0x15, 0x24, 0x1E, 0x6D, 0x5D, 0x51, 0x0A, 0x2D, 0x75, 0x38, 0x26, 0x56,
	0x1B, 0x1A, 0x1C, 0x03, 0x5C, 0x3C, 0x28, 0x0D, 0x38, 0x04, 0x40, 0x1B,
	0x2D, 0x17, 0x1E, 0x00, 0x15, 0x3A, 0x18, 0x36, 0x29, 0x0A, 0x07, 0x17,
	0x08, 0x5F, 0x16, 0x0D, 0x3B, 0x20, 0x59, 0x71, 0x09, 0x27, 0x22, 0x12,
	0x2E, 0x3C, 0x03, 0x1F, 0x1F, 0x74, 0x16, 0x54, 0x22, 0x1E, 0x30, 0x3F,
	0x26, 0x0B, 0x52, 0x08, 0x20, 0x03, 0x29, 0x5C, 0x2E, 0x0E, 0x30, 0x3D,
	0x1A, 0x74, 0x54, 0x03, 0x16, 0x2F, 0x16, 0x24, 0x36, 0x25, 0x53, 0x15,
	0x59, 0x03, 0x36, 0x0D, 0x0B, 0x16, 0x52, 0x5E, 0x1F, 0x73, 0x54, 0x35,
	0x41, 0x0D, 0x74, 0x19, 0x05, 0x07, 0x06, 0x2D, 0x28, 0x02, 0x37, 0x3F,
	0x74, 0x39, 0x16, 0x25, 0x53, 0x12, 0x3F, 0x4E, 0x27, 0x33, 0x30, 0x03,
	0x05, 0x28, 0x08, 0x2F, 0x5C, 0x26, 0x08, 0x53, 0x0D, 0x3C, 0x50, 0x38,
	0x58, 0x75, 0x23, 0x2F, 0x06, 0x24, 0x2D, 0x5F, 0x00, 0x39, 0x24, 0x07,
	0x5C, 0x36, 0x0D, 0x24, 0x32, 0x25, 0x04, 0x1B, 0x25, 0x76, 0x18, 0x50,
	0x3E, 0x3F, 0x29, 0x36, 0x18, 0x22, 0x3D, 0x12, 0x3A, 0x2D, 0x5E, 0x20,
	0x31, 0x29, 0x22, 0x36, 0x05, 0x26, 0x25, 0x23, 0x3A, 0x0D, 0x74, 0x1A,
	0x34, 0x3A, 0x2E, 0x77, 0x5C, 0x27, 0x2A, 0x0F, 0x32, 0x5C, 0x09, 0x2A,
	0x27, 0x16, 0x07, 0x2C, 0x0A, 0x0F, 0x13, 0x19, 0x37, 0x07, 0x2D, 0x24,
	0x15, 0x00, 0x29, 0x53, 0x26, 0x00, 0x10, 0x39, 0x5B, 0x33, 0x5D, 0x29,
	0x00, 0x0A, 0x00, 0x36, 0x22, 0x2F, 0x2D, 0x2F, 0x3A, 0x03, 0x0D, 0x2A,
	0x18, 0x1F, 0x22, 0x06, 0x2D, 0x0E, 0x35, 0x27, 0x3B, 0x0E, 0x33, 0x3F,
	0x57, 0x3C, 0x28, 0x20, 0x1C, 0x52, 0x23, 0x04, 0x07, 0x1F, 0x50, 0x5D,
	0x00, 0x16, 0x3A, 0x18, 0x01, 0x5A, 0x2A, 0x5D, 0x0F, 0x0C, 0x5C, 0x30,
	0x3B, 0x35, 0x19, 0x25, 0x70, 0x21, 0x24, 0x1D, 0x24, 0x27, 0x3D, 0x53,
	0x03, 0x26, 0x2E, 0x47, 0x2D, 0x01, 0x0F, 0x35, 0x06, 0x52, 0x25, 0x31,
	0x24, 0x5F, 0x34, 0x38, 0x3F, 0x29, 0x47, 0x05, 0x07, 0x0C, 0x0F, 0x39,
	0x4A, 0x3D, 0x1B, 0x74, 0x08, 0x12, 0x2F, 0x33, 0x03, 0x43, 0x28, 0x21,
	0x22, 0x26, 0x2F, 0x0C, 0x0B, 0x3A, 0x7A, 0x25, 0x57, 0x0C, 0x18, 0x26,
	0x5A, 0x29, 0x26, 0x1C, 0x05, 0x2B, 0x55, 0x01, 0x27, 0x34, 0x3C, 0x53,
	0x3F, 0x03, 0x12, 0x0B, 0x11, 0x24, 0x2D, 0x1B, 0x3E, 0x06, 0x5B, 0x3C,
	0x75, 0x1F, 0x02, 0x21, 0x0D, 0x09, 0x22, 0x32, 0x02, 0x32, 0x76, 0x16,
	0x16, 0x39, 0x05, 0x2B, 0x47, 0x57, 0x1A, 0x31, 0x6D, 0x55, 0x19, 0x39,
	0x3B, 0x2F, 0x38, 0x04, 0x20, 0x21, 0x2E, 0x26, 0x29, 0x1B, 0x01, 0x00,
	0x14, 0x54, 0x25, 0x28, 0x23, 0x1E, 0x10, 0x5D, 0x0F, 0x71, 0x28, 0x3B,
	0x1A, 0x2F, 0x23, 0x3A, 0x38, 0x1B, 0x20, 0x69, 0x06, 0x33, 0x0D, 0x06,
	0x23, 0x22, 0x3B, 0x09, 0x3D, 0x77, 0x18, 0x34, 0x1D, 0x04, 0x72, 0x3F,
	0x2C, 0x2D, 0x32, 0x29, 0x21, 0x2E, 0x41, 0x18, 0x04, 0x29, 0x25, 0x24,
	0x03, 0x3A, 0x38, 0x2A, 0x5D, 0x59, 0x36, 0x38, 0x28, 0x3D, 0x20, 0x37,
	0x1D, 0x37, 0x02, 0x1B, 0x04, 0x54, 0x0E, 0x2A, 0x05, 0x12, 0x2D, 0x12,
	0x17, 0x2A, 0x21, 0x16, 0x22, 0x3A, 0x1E, 0x2C, 0x1A, 0x28, 0x5B, 0x02,
	0x23, 0x2B, 0x09, 0x08, 0x28, 0x21, 0x25, 0x0E, 0x5C, 0x21, 0x0A, 0x19,
	0x35, 0x29, 0x40, 0x24, 0x3F, 0x0D, 0x24, 0x06, 0x73, 0x39, 0x24, 0x25,
	0x59, 0x74, 0x35, 0x07, 0x37, 0x18, 0x26, 0x08, 0x55, 0x5C, 0x2A, 0x31,
	0x21, 0x51, 0x22, 0x19, 0x16, 0x39, 0x11, 0x38, 0x2C, 0x32, 0x35, 0x23,
	0x3E, 0x18, 0x33, 0x3F, 0x0E, 0x2B, 0x0C, 0x12, 0x0A, 0x10, 0x00, 0x3D,
	0x7B, 0x38, 0x29, 0x5D, 0x00, 0x09, 0x3B, 0x06, 0x56, 0x26, 0x77, 0x23,
	0x24, 0x1F, 0x1D, 0x13, 0x5C, 0x33, 0x16, 0x3E, 0x77, 0x01, 0x1B, 0x5E,
	0x27, 0x31, 0x2F, 0x36, 0x2D, 0x27, 0x11, 0x5B, 0x0B, 0x45, 0x06, 0x23,
	0x02, 0x39, 0x0F, 0x38, 0x10, 0x03, 0x34, 0x06, 0x2F, 0x3A, 0x5D, 0x31,
	0x39, 0x2E, 0x74, 0x05, 0x2F, 0x45, 0x0F, 0x21, 0x39, 0x58, 0x25, 0x59,
	0x2D, 0x29, 0x33, 0x39, 0x5E, 0x2E, 0x1B, 0x26, 0x2F, 0x52, 0x32, 0x00,
	0x53, 0x04, 0x26, 0x2C, 0x2F, 0x27, 0x19, 0x20, 0x76, 0x2A, 0x2D, 0x1A,
	0x28, 0x13, 0x36, 0x18, 0x2F, 0x0E, 0x10, 0x1D, 0x0B, 0x14, 0x2E, 0x35,
	0x2B, 0x12, 0x2C, 0x04, 0x30, 0x36, 0x32, 0x2C, 0x02, 0x35, 0x2E, 0x02,
	0x1E, 0x21, 0x17, 0x1B, 0x02, 0x2D, 0x2C, 0x03, 0x2F, 0x56, 0x38, 0x09,
	0x05, 0x3E, 0x06, 0x21, 0x32, 0x0E, 0x06, 0x0C, 0x21, 0x18, 0x07, 0x5A,
	0x51, 0x20, 0x3B, 0x24, 0x03, 0x32, 0x59, 0x5F, 0x11, 0x54, 0x26, 0x2C,
	0x5A, 0x31, 0x14, 0x55, 0x0F, 0x23, 0x1B, 0x59, 0x4A, 0x34, 0x5A, 0x16,
	0x5F, 0x59, 0x1D, 0x00, 0x75, 0x0A, 0x04, 0x0C, 0x29, 0x06, 0x2F, 0x51,
	0x2B, 0x13, 0x14, 0x3D, 0x24, 0x26, 0x1E, 0x1A, 0x58, 0x38, 0x3C, 0x12,
	0x0C, 0x3D, 0x0A, 0x59, 0x31, 0x09, 0x16, 0x54, 0x39, 0x22, 0x08, 0x05,
	0x2F, 0x14, 0x26, 0x33, 0x0B, 0x32, 0x3A, 0x3E, 0x70, 0x5F, 0x59, 0x03,
	0x00, 0x06, 0x1A, 0x34, 0x5C, 0x0F, 0x13, 0x2D, 0x32, 0x27, 0x04, 0x11,
	0x5D, 0x20, 0x5C, 0x52, 0x1A, 0x19, 0x54, 0x39, 0x19, 0x74, 0x23, 0x39,
	0x29, 0x2A, 0x31, 0x35, 0x11, 0x02, 0x03, 0x24, 0x3E, 0x00, 0x28, 0x11,
	0x08, 0x1F, 0x50, 0x57, 0x40, 0x37, 0x0E, 0x03, 0x20, 0x1F, 0x33, 0x07,
	0x38, 0x21, 0x1F, 0x34, 0x1D, 0x08, 0x2D, 0x1E, 0x05, 0x34, 0x27, 0x07,
	0x1C, 0x12, 0x1D, 0x03, 0x39, 0x12, 0x29, 0x58, 0x33, 0x5F, 0x5B, 0x7B,
	0x1E, 0x50, 0x26, 0x1B, 0x21, 0x1D, 0x23, 0x5E, 0x24, 0x26, 0x1C, 0x58,
	0x16, 0x1C, 0x29, 0x21, 0x23, 0x3A, 0x29, 0x17, 0x19, 0x54, 0x21, 0x29,
	0x26, 0x2D, 0x25, 0x1E, 0x59, 0x31, 0x5C, 0x2C, 0x1E, 0x2A, 0x00, 0x25,
	0x51, 0x34, 0x1C, 0x0F, 0x5C, 0x31, 0x16, 0x3C, 0x69, 0x43, 0x0D, 0x16,
	0x2C, 0x25, 0x29, 0x18, 0x18, 0x58, 0x7A, 0x21, 0x0D, 0x0A, 0x18, 0x69,
	0x5C, 0x19, 0x08, 0x5B, 0x69, 0x54, 0x0A, 0x0B, 0x40, 0x0C, 0x54, 0x26,
	0x17, 0x06, 0x76, 0x2D, 0x39, 0x07, 0x5C, 0x26, 0x00, 0x18, 0x37, 0x24,
	0x12, 0x3D, 0x26, 0x1F, 0x53, 0x12, 0x26, 0x0C, 0x3E, 0x2D, 0x37, 0x15,
	0x26, 0x14, 0x3F, 0x28, 0x59, 0x32, 0x0B, 0x5A, 0x34, 0x0B, 0x08, 0x02,
	0x22, 0x29, 0x25, 0x10, 0x01, 0x05, 0x23, 0x0F, 0x06, 0x3F, 0x1C, 0x03,
	0x2B, 0x05, 0x1C, 0x33, 0x07, 0x36, 0x10, 0x0B, 0x0A, 0x2C, 0x5C, 0x10,
	0x00, 0x1E, 0x27, 0x3B, 0x57, 0x1F, 0x26, 0x0A, 0x2E, 0x12, 0x56, 0x02,
	0x01, 0x47, 0x13, 0x56, 0x5A, 0x2B, 0x3A, 0x52, 0x3D, 0x31, 0x17, 0x55,
	0x04, 0x2D, 0x19, 0x6D, 0x03, 0x07, 0x29, 0x0C, 0x25, 0x59, 0x04, 0x27,
	0x20, 0x3B, 0x54, 0x32, 0x0A, 0x26, 0x21, 0x2D, 0x24, 0x27, 0x5E, 0x69,
	0x38, 0x33, 0x5A, 0x3E, 0x7A, 0x1B, 0x2D, 0x19, 0x38, 0x05, 0x59, 0x2F,
	0x00, 0x0C, 0x2E, 0x58, 0x20, 0x56, 0x32, 0x2F, 0x3D, 0x2E, 0x14, 0x04,
	0x24, 0x06, 0x2A, 0x3D, 0x1B, 0x28, 0x2A, 0x32, 0x57, 0x29, 0x28, 0x16,
	0x55, 0x20, 0x0F, 0x07, 0x3F, 0x06, 0x5B, 0x01, 0x29, 0x28, 0x33, 0x0A,
	0x1F, 0x77, 0x19, 0x12, 0x04, 0x11, 0x75, 0x09, 0x17, 0x26, 0x5D, 0x77,
	0x07, 0x0A, 0x14, 0x0D, 0x21, 0x1B, 0x20, 0x3B, 0x33, 0x6D, 0x00, 0x24,
	0x34, 0x31, 0x7A, 0x34, 0x17, 0x39, 0x1D, 0x35, 0x35, 0x37, 0x3E, 0x5B,
	0x3A, 0x3F, 0x34, 0x5D, 0x2F, 0x25, 0x09, 0x37, 0x1D, 0x01, 0x74, 0x38,
	0x16, 0x1C, 0x08, 0x34, 0x0A, 0x30, 0x59, 0x22, 0x30, 0x02, 0x4E, 0x2B,
	0x0D, 0x0A, 0x25, 0x2E, 0x27, 0x5A, 0x31, 0x0E, 0x24, 0x2A, 0x0F, 0x01,
	0x05, 0x0A, 0x3E, 0x22, 0x38, 0x1E, 0x34, 0x0B, 0x31, 0x0F, 0x43, 0x02,
	0x34, 0x3A, 0x17, 0x00, 0x20, 0x1C, 0x1B, 0x27, 0x16, 0x24, 0x21, 0x1D,
	0x30, 0x15, 0x37, 0x41, 0x40, 0x6D, 0x0A, 0x26, 0x0D, 0x2C, 0x20, 0x55,
	0x34, 0x2C, 0x31, 0x18, 0x55, 0x2C, 0x59, 0x3C, 0x1A, 0x3A, 0x27, 0x45,
	0x20, 0x3A, 0x1A, 0x29, 0x1A, 0x01, 0x3B, 0x3E, 0x0A, 0x23, 0x28, 0x35,
	0x26, 0x08, 0x1E, 0x44, 0x0C, 0x20, 0x25, 0x5A, 0x13, 0x0F, 0x1D, 0x19,
	0x07, 0x38, 0x2F, 0x0E, 0x0C, 0x41, 0x19, 0x7B, 0x5B, 0x05, 0x0A, 0x23,
	0x34, 0x5F, 0x50, 0x3F, 0x24, 0x36, 0x54, 0x16, 0x5A, 0x26, 0x37, 0x28,
	0x4A, 0x57, 0x52, 0x06, 0x25, 0x03, 0x5E, 0x52, 0x74, 0x3A, 0x33, 0x2D,
	0x2A, 0x24, 0x22, 0x25, 0x06, 0x38, 0x1B, 0x5F, 0x2D, 0x06, 0x02, 0x17,
	0x5C, 0x0E, 0x3A, 0x40, 0x09, 0x3E, 0x2E, 0x3E, 0x03, 0x37, 0x14, 0x20,
	0x02, 0x11, 0x2A, 0x1E, 0x27, 0x07, 0x38, 0x3A, 0x09, 0x06, 0x27, 0x3D,
	0x7A, 0x1A, 0x27, 0x0C, 0x32, 0x01, 0x14, 0x58, 0x45, 0x07, 0x6D, 0x07,
	0x2E, 0x45, 0x05, 0x1B, 0x1A, 0x53, 0x03, 0x5C, 0x24, 0x15, 0x58, 0x14,
	0x3E, 0x0D, 0x01, 0x18, 0x1B, 0x29, 0x14, 0x06, 0x51, 0x25, 0x3D, 0x75,
	0x3A, 0x1B, 0x5B, 0x21, 0x03, 0x05, 0x16, 0x0A, 0x3B, 0x14, 0x21, 0x36,
	0x17, 0x3C, 0x2E, 0x14, 0x23, 0x57, 0x19, 0x16, 0x5B, 0x29, 0x07, 0x2C,
	0x30, 0x3C, 0x58, 0x19, 0x3A, 0x14, 0x3C, 0x02, 0x08, 0x06, 0x00, 0x3F,
	0x29, 0x07, 0x3F, 0x09, 0x5F, 0x24, 0x5C, 0x3C, 0x2C, 0x27, 0x04, 0x59,
	0x1B, 0x2E, 0x1B, 0x0F, 0x45, 0x3E, 0x70, 0x0E, 0x4E, 0x01, 0x3E, 0x38,
	0x22, 0x2E, 0x0F, 0x0F, 0x0F, 0x0B, 0x08, 0x1E, 0x1A, 0x03, 0x54, 0x31,
	0x3C, 0x40, 0x69, 0x39, 0x54, 0x19, 0x58, 0x35, 0x38, 0x24, 0x02, 0x05,
	0x34, 0x5F, 0x39, 0x3E, 0x07, 0x0D, 0x47, 0x05, 0x59, 0x31, 0x2F, 0x15,
	0x25, 0x2A, 0x5A, 0x16, 0x24, 0x0B, 0x38, 0x28, 0x23, 0x00, 0x2C, 0x19,
	0x12, 0x7A, 0x2B, 0x25, 0x3C, 0x1E, 0x20, 0x19, 0x33, 0x14, 0x5C, 0x37,
	0x34, 0x1B, 0x34, 0x2D, 0x75, 0x3B, 0x55, 0x5C, 0x2C, 0x05, 0x25, 0x4A,
	0x25, 0x09, 0x0D, 0x2A, 0x33, 0x24, 0x40, 0x17, 0x18, 0x06, 0x06, 0x2E,
	0x69, 0x0A, 0x14, 0x0C, 0x1E, 0x05, 0x3A, 0x38, 0x0F, 0x1A, 0x69, 0x23,
	0x0D, 0x1D, 0x5A, 0x73, 0x1B, 0x19, 0x3C, 0x12, 0x25, 0x2A, 0x17, 0x25,
	0x11, 0x14, 0x0F, 0x18, 0x1A, 0x5E, 0x16, 0x38, 0x55, 0x45, 0x3E, 0x35,
	0x1C, 0x34, 0x21, 0x2C, 0x6D, 0x3B, 0x03, 0x5E, 0x5D, 0x76, 0x0E, 0x0F,
	0x28, 0x25, 0x1A, 0x18, 0x54, 0x41, 0x0E, 0x75, 0x1C, 0x0F, 0x14, 0x12,
	0x0A, 0x1E, 0x2D, 0x0C, 0x59, 0x21, 0x23, 0x2C, 0x20, 0x2C, 0x72, 0x1A,
	0x19, 0x59, 0x13, 0x16, 0x05, 0x0D, 0x3B, 0x1D, 0x17, 0x22, 0x18, 0x0D,
	0x22, 0x69, 0x3F, 0x09, 0x5B, 0x58, 0x74, 0x0A, 0x53, 0x5F, 0x44, 0x25,
	0x54, 0x18, 0x0B, 0x03, 0x29, 0x54, 0x10, 0x05, 0x39, 0x03, 0x09, 0x37,
	0x25, 0x13, 0x17, 0x07, 0x30, 0x19, 0x40, 0x17, 0x2B, 0x52, 0x36, 0x11,
	0x33, 0x21, 0x07, 0x39, 0x00, 0x6D, 0x54, 0x2B, 0x21, 0x00, 0x77, 0x3B,
	0x15, 0x02, 0x0C, 0x35, 0x18, 0x23, 0x3A, 0x3E, 0x0F, 0x06, 0x17, 0x17,
	0x0C, 0x2A, 0x1E, 0x28, 0x17, 0x1B, 0x21, 0x3C, 0x38, 0x5D, 0x21, 0x38,
	0x34, 0x16, 0x3B, 0x22, 0x7A, 0x18, 0x17, 0x5E, 0x06, 0x7A, 0x39, 0x28,
	0x2D, 0x40, 0x30, 0x04, 0x1B, 0x0D, 0x21, 0x0A, 0x5A, 0x23, 0x28, 0x38,
	0x17, 0x29, 0x13, 0x1E, 0x1E, 0x0F, 0x39, 0x15, 0x20, 0x0A, 0x2D, 0x22,
	0x23, 0x07, 0x31, 0x70, 0x21, 0x38, 0x18, 0x00, 0x32, 0x5D, 0x25, 0x5F,
	0x11, 0x74, 0x0A, 0x0B, 0x0A, 0x02, 0x16, 0x15, 0x29, 0x1C, 0x3E, 0x72,
	0x01, 0x07, 0x25, 0x19, 0x38, 0x39, 0x0E, 0x5A, 0x33, 0x69, 0x22, 0x32,
	0x0F, 0x0C, 0x35, 0x2E, 0x31, 0x21, 0x05, 0x14, 0x29, 0x37, 0x28, 0x1F,
	0x0B, 0x55, 0x0B, 0x59, 0x59, 0x3B, 0x07, 0x27, 0x3B, 0x13, 0x23, 0x39,
	0x19, 0x3B, 0x44, 0x27, 0x20, 0x56, 0x18, 0x39, 0x1A, 0x09, 0x00, 0x41,
	0x0D, 0x25, 0x43, 0x25, 0x56, 0x5A, 0x0A, 0x01, 0x26, 0x18, 0x44, 0x17,
	0x3B, 0x4E, 0x2F, 0x1A, 0x06, 0x0F, 0x15, 0x16, 0x29, 0x20, 0x59, 0x57,
	0x2C, 0x07, 0x74, 0x1C, 0x2D, 0x5B, 0x5B, 0x0A, 0x5B, 0x52, 0x3E, 0x3B,
	0x17, 0x0D, 0x16, 0x41, 0x27, 0x27, 0x27, 0x2D, 0x02, 0x3F, 0x33, 0x1B,
	0x36, 0x28, 0x3C, 0x0E, 0x58, 0x12, 0x38, 0x38, 0x76, 0x25, 0x53, 0x39,
	0x38, 0x7B, 0x47, 0x07, 0x1A, 0x3B, 0x7A, 0x22, 0x04, 0x20, 0x5E, 0x77,
	0x36, 0x0E, 0x2D, 0x5C, 0x38, 0x36, 0x10, 0x37, 0x5E, 0x6D, 0x0B, 0x15,
	0x28, 0x31, 0x08, 0x0A, 0x59, 0x2C, 0x1E, 0x17, 0x01, 0x15, 0x5B, 0x04,
	0x71, 0x43, 0x17, 0x0B, 0x01, 0x36, 0x22, 0x08, 0x02, 0x3A, 0x23, 0x1A,
	0x11, 0x5B, 0x32, 0x31, 0x1A, 0x35, 0x56, 0x18, 0x14, 0x02, 0x52, 0x24,
	0x2C, 0x31, 0x3C, 0x1B, 0x0D, 0x26, 0x3A, 0x2F, 0x07, 0x5C, 0x19, 0x27,
	0x25, 0x0C, 0x0C, 0x0C, 0x18, 0x55, 0x29, 0x20, 0x02, 0x2C, 0x24, 0x0F,
	0x2C, 0x2A, 0x70, 0x2A, 0x05, 0x08, 0x18, 0x6D, 0x5A, 0x18, 0x22, 0x0F,
	0x05, 0x2A, 0x58, 0x2D, 0x38, 0x3B, 0x3F, 0x18, 0x5C, 0x3E, 0x26, 0x38,
	0x13, 0x5B, 0x3D, 0x7B, 0x04, 0x0D, 0x27, 0x12, 0x0C, 0x3D, 0x3B, 0x19,
	0x25, 0x3B, 0x07, 0x11, 0x34, 0x2E, 0x1A, 0x0F, 0x4A, 0x1E, 0x5D, 0x00,
	0x0A, 0x26, 0x0A, 0x32, 0x21, 0x2F, 0x37, 0x16, 0x1D, 0x0B, 0x38, 0x39,
	0x5F, 0x01, 0x73, 0x2B, 0x57, 0x1D, 0x2C, 0x7B, 0x0B, 0x0D, 0x3F, 0x38,
	0x26, 0x36, 0x37, 0x56, 0x01, 0x32, 0x3B, 0x2F, 0x28, 0x5D, 0x06, 0x0B,
	0x15, 0x04, 0x3E, 0x27, 0x20, 0x53, 0x57, 0x2C, 0x36, 0x59, 0x00, 0x28,
	0x2E, 0x35, 0x3A, 0x25, 0x1D, 0x44, 0x05, 0x5A, 0x30, 0x3F, 0x33, 0x14,
	0x34, 0x18, 0x45, 0x44, 0x29, 0x1E, 0x35, 0x27, 0x0A, 0x07, 0x5A, 0x17,
	0x01, 0x25, 0x31, 0x2D, 0x0F, 0x5C, 0x33, 0x6D, 0x23, 0x53, 0x29, 0x2A,
	0x6D, 0x3F, 0x58, 0x34, 0x23, 0x37, 0x21, 0x05, 0x34, 0x3B, 0x21, 0x26,
	0x23, 0x18, 0x33, 0x34, 0x5F, 0x34, 0x19, 0x26, 0x0A, 0x27, 0x54, 0x09,
	0x13, 0x28, 0x3A, 0x51, 0x1C, 0x04, 0x21, 0x54, 0x53, 0x57, 0x2A, 0x13,
	0x1C, 0x07, 0x0F, 0x08, 0x73, 0x04, 0x52, 0x37, 0x38, 0x2C, 0x27, 0x35,
	0x38, 0x2D, 0x69, 0x5A, 0x3B, 0x23, 0x2C, 0x2B, 0x1F, 0x0E, 0x39, 0x27,
	0x3A, 0x07, 0x15, 0x17, 0x08, 0x31, 0x1A, 0x51, 0x1A, 0x29, 0x36, 0x08,
	0x03, 0x03, 0x1D, 0x38, 0x55, 0x28, 0x16, 0x29, 0x72, 0x36, 0x1B, 0x26,
	0x59, 0x23, 0x0A, 0x11, 0x29, 0x19, 0x7A, 0x55, 0x59, 0x0B, 0x44, 0x27,
	0x38, 0x58, 0x57, 0x1F, 0x2E, 0x03, 0x30, 0x03, 0x1A, 0x24, 0x1E, 0x34,
	0x5A, 0x13, 0x70, 0x08, 0x2A, 0x56, 0x53, 0x36, 0x38, 0x50, 0x19, 0x21,
	0x7A, 0x1D, 0x30, 0x27, 0x0A, 0x2C, 0x1E, 0x26, 0x3E, 0x5B, 0x2F, 0x09,
	0x17, 0x3E, 0x03, 0x05, 0x03, 0x0B, 0x16, 0x21, 0x16, 0x14, 0x30, 0x00,
	0x33, 0x35, 0x54, 0x34, 0x24, 0x11, 0x7A, 0x00, 0x33, 0x59, 0x3F, 0x1A,
	0x16, 0x54, 0x27, 0x01, 0x0E, 0x1B, 0x23, 0x1C, 0x27, 0x12, 0x00, 0x0F,
	0x18, 0x13, 0x38, 0x59, 0x2E, 0x56, 0x1A, 0x10, 0x1A, 0x2E, 0x17, 0x11,
	0x77, 0x39, 0x0B, 0x1A, 0x0D, 0x3B, 0x18, 0x29, 0x18, 0x1D, 0x31, 0x02,
	0x0A, 0x17, 0x25, 0x2D, 0x2F, 0x29, 0x09, 0x08, 0x1A, 0x36, 0x0F, 0x41,
	0x1E, 0x75, 0x2A, 0x07, 0x07, 0x20, 0x11, 0x09, 0x2D, 0x3B, 0x3F, 0x37,
	0x0A, 0x0B, 0x5E, 0x1E, 0x10, 0x2B, 0x55, 0x5B, 0x38, 0x76, 0x0B, 0x59,
	0x0A, 0x2F, 0x29, 0x38, 0x28, 0x1A, 0x0D, 0x0D, 0x3D, 0x4A, 0x59, 0x0E,
	0x7B, 0x02, 0x11, 0x23, 0x0D, 0x37, 0x2D, 0x05, 0x09, 0x24, 0x2D, 0x38,
	0x16, 0x16, 0x27, 0x29, 0x14, 0x18, 0x5F, 0x26, 0x24, 0x19, 0x32, 0x5F,
	0x1A, 0x3B, 0x0A, 0x4E, 0x5D, 0x28, 0x7A, 0x54, 0x0C, 0x2D, 0x2D, 0x13,
	0x38, 0x15, 0x5C, 0x09, 0x12, 0x15, 0x51, 0x56, 0x20, 0x2F, 0x20, 0x22,
	0x27, 0x58, 0x2B, 0x23, 0x39, 0x00, 0x09, 0x34, 0x0A, 0x39, 0x19, 0x1D,
	0x37, 0x47, 0x52, 0x2C, 0x2A, 0x20, 0x5D, 0x12, 0x5D, 0x23, 0x71, 0x14,
	0x39, 0x00, 0x09, 0x2E, 0x0B, 0x53, 0x0D, 0x27, 0x28, 0x59, 0x31, 0x18,
	0x53, 0x0F, 0x20, 0x0B, 0x22, 0x03, 0x00, 0x43, 0x2F, 0x0D, 0x01, 0x09,
	0x07, 0x57, 0x20, 0x52, 0x08, 0x2E, 0x05, 0x1B, 0x3A, 0x72, 0x19, 0x30,
	0x2C, 0x23, 0x2E, 0x04, 0x2E, 0x27, 0x44, 0x08, 0x05, 0x4E, 0x02, 0x26,
	0x1A, 0x19, 0x18, 0x18, 0x02, 0x7A, 0x01, 0x2D, 0x20, 0x22, 0x3B, 0x47,
	0x30, 0x09, 0x2D, 0x77, 0x5C, 0x2C, 0x08, 0x00, 0x10, 0x34, 0x2F, 0x0A,
	0x3F, 0x04, 0x5B, 0x06, 0x1E, 0x32, 0x1A, 0x1D, 0x17, 0x08, 0x29, 0x09,
	0x34, 0x35, 0x27, 0x3E, 0x71, 0x07, 0x59, 0x5B, 0x07, 0x75, 0x16, 0x55,
	0x22, 0x3D, 0x69, 0x3F, 0x2B, 0x56, 0x18, 0x0A, 0x00, 0x26, 0x3A, 0x3C,
	0x20, 0x47, 0x2C, 0x02, 0x06, 0x13, 0x18, 0x17, 0x17, 0x26, 0x17, 0x1E,
	0x59, 0x23, 0x59, 0x20, 0x1E, 0x59, 0x28, 0x11, 0x08, 0x15, 0x02, 0x18,
	0x40, 0x34, 0x02, 0x39, 0x5F, 0x53, 0x69, 0x43, 0x17, 0x04, 0x5E, 0x2D,
	0x04, 0x13, 0x27, 0x5C, 0x1B, 0x04, 0x19, 0x56, 0x23, 0x7B, 0x3E, 0x58,
	0x5F, 0x3C, 0x34, 0x29, 0x16, 0x38, 0x52, 0x31, 0x47, 0x31, 0x2B, 0x39,
	0x0F, 0x3A, 0x52, 0x5A, 0x12, 0x10, 0x24, 0x33, 0x5F, 0x53, 0x6D, 0x26,
	0x04, 0x29, 0x5E, 0x31, 0x5E, 0x50, 0x03, 0x03, 0x0F, 0x0A, 0x54, 0x21,
	0x0D, 0x76, 0x5F, 0x0F, 0x0C, 0x52, 0x0A, 0x5B, 0x22, 0x25, 0x1D, 0x01,
	0x22, 0x00, 0x41, 0x5A, 0x7A, 0x16, 0x08, 0x58, 0x3D, 0x2E, 0x27, 0x2D,
	0x1D, 0x1D, 0x76, 0x1A, 0x04, 0x20, 0x12, 0x7A, 0x58, 0x04, 0x17, 0x13,
	0x7A, 0x03, 0x31, 0x5D, 0x40, 0x7B, 0x01, 0x02, 0x38, 0x3B, 0x2F, 0x2E,
	0x03, 0x3E, 0x5C, 0x1B, 0x3C, 0x4A, 0x24, 0x18, 0x24, 0x1A, 0x2F, 0x34,
	0x09, 0x04, 0x58, 0x1B, 0x00, 0x19, 0x0A, 0x59, 0x1B, 0x56, 0x06, 0x24,
	0x1E, 0x0C, 0x00, 0x44, 0x12, 0x14, 0x08, 0x08, 0x07, 0x3B, 0x55, 0x35,
	0x41, 0x59, 0x32, 0x23, 0x55, 0x26, 0x2C, 0x74, 0x00, 0x25, 0x23, 0x59,
	0x10, 0x01, 0x00, 0x56, 0x2E, 0x12, 0x0A, 0x06, 0x59, 0x22, 0x10, 0x1D,
	0x4E, 0x18, 0x28, 0x24, 0x14, 0x2E, 0x27, 0x5A, 0x35, 0x23, 0x28, 0x5F,
	0x5E, 0x70, 0x28, 0x19, 0x38, 0x0E, 0x25, 0x2D, 0x2A, 0x37, 0x23, 0x04,
	0x29, 0x08, 0x1E, 0x3A, 0x15, 0x16, 0x14, 0x23, 0x52, 0x07, 0x0A, 0x06,
	0x16, 0x5A, 0x26, 0x43, 0x28, 0x26, 0x5C, 0x31, 0x0A, 0x20, 0x3E, 0x23,
	0x35, 0x34, 0x4E, 0x29, 0x06, 0x0D, 0x58, 0x09, 0x34, 0x27, 0x32, 0x21,
	0x31, 0x14, 0x2F, 0x14, 0x43, 0x00, 0x19, 0x12, 0x20, 0x43, 0x54, 0x00,
	0x01, 0x0D, 0x02, 0x4A, 0x09, 0x5B, 0x3A, 0x5F, 0x55, 0x09, 0x05, 0x76,
	0x0F, 0x51, 0x0F, 0x2E, 0x7B, 0x5A, 0x4E, 0x28, 0x06, 0x13, 0x58, 0x54,
	0x18, 0x5E, 0x6D, 0x14, 0x07, 0x04, 0x31, 0x24, 0x36, 0x1B, 0x21, 0x07,
	0x33, 0x29, 0x2D, 0x00, 0x1D, 0x0E, 0x00, 0x2D, 0x2B, 0x05, 0x29, 0x3E,
	0x0C, 0x0B, 0x40, 0x7A, 0x47, 0x39, 0x26, 0x06, 0x0F, 0x15, 0x19, 0x02,
	0x58, 0x17, 0x04, 0x58, 0x1B, 0x13, 0x75, 0x5A, 0x1B, 0x07, 0x5B, 0x69,
	0x15, 0x37, 0x57, 0x3E, 0x2D, 0x3A, 0x56, 0x45, 0x23, 0x16, 0x3A, 0x18,
	0x22, 0x04, 0x25, 0x03, 0x03, 0x38, 0x19, 0x24, 0x2D, 0x26, 0x34, 0x2E,
	0x0D, 0x34, 0x50, 0x1B, 0x0D, 0x36, 0x1B, 0x14, 0x2A, 0x21, 0x11, 0x02,
	0x11, 0x5F, 0x5F, 0x2E, 0x0E, 0x13, 0x14, 0x1B, 0x0A, 0x43, 0x59, 0x3E,
	0x5E, 0x01, 0x01, 0x2C, 0x27, 0x28, 0x06, 0x21, 0x24, 0x07, 0x1B, 0x31,
	0x3C, 0x19, 0x5B, 0x1D, 0x25, 0x0D, 0x16, 0x56, 0x52, 0x69, 0x03, 0x54,
	0x5B, 0x0E, 0x2F, 0x35, 0x17, 0x41, 0x0D, 0x38, 0x5E, 0x0C, 0x36, 0x22,
	0x23, 0x43, 0x14, 0x26, 0x05, 0x0F, 0x5D, 0x13, 0x22, 0x44, 0x3B, 0x5F,
	0x17, 0x22, 0x09, 0x69, 0x5B, 0x54, 0x19, 0x53, 0x0E, 0x34, 0x0C, 0x5D,
	0x05, 0x7B, 0x24, 0x4A, 0x0A, 0x01, 0x23, 0x06, 0x3B, 0x0C, 0x53, 0x23,
	0x36, 0x56, 0x3D, 0x02, 0x31, 0x14, 0x0B, 0x1A, 0x5B, 0x29, 0x1F, 0x38,
	0x01, 0x44, 0x70, 0x21, 0x54, 0x21, 0x05, 0x06, 0x1E, 0x4A, 0x1E, 0x53,
	0x14, 0x1D, 0x11, 0x0B, 0x25, 0x3B, 0x3F, 0x23, 0x14, 0x5B, 0x76, 0x35,
	0x38, 0x1C, 0x27, 0x72, 0x0E, 0x59, 0x41, 0x2D, 0x2F, 0x09, 0x19, 0x58,
	0x33, 0x0E, 0x0A, 0x00, 0x56, 0x25, 0x0C, 0x21, 0x50, 0x04, 0x5D, 0x13,
	0x15, 0x05, 0x3A, 0x21, 0x15, 0x39, 0x18, 0x21, 0x09, 0x27, 0x03, 0x0B,
	0x18, 0x40, 0x0D, 0x1D, 0x50, 0x23, 0x1D, 0x76, 0x5A, 0x18, 0x5D, 0x5F,
	0x27, 0x21, 0x38, 0x29, 0x13, 0x2E, 0x43, 0x0D, 0x36, 0x1D, 0x14, 0x22,
	0x29, 0x14, 0x19, 0x2C, 0x35, 0x13, 0x14, 0x5A, 0x6D, 0x3B, 0x12, 0x16,
	0x58, 0x36, 0x1D, 0x2A, 0x18, 0x3B, 0x17, 0x5C, 0x17, 0x28, 0x27, 0x6D,
	0x07, 0x06, 0x00, 0x1D, 0x71, 0x43, 0x0A, 0x3C, 0x58, 0x34, 0x1E, 0x0C,
	0x00, 0x19, 0x0C, 0x58, 0x10, 0x58, 0x2C, 0x17, 0x59, 0x57, 0x5F, 0x25,
	0x7B, 0x54, 0x33, 0x5B, 0x0A, 0x71, 0x5E, 0x11, 0x14, 0x07, 0x37, 0x5F,
	0x03, 0x45, 0x11, 0x2C, 0x1E, 0x38, 0x45, 0x3B, 0x07, 0x5E, 0x4A, 0x5F,
	0x44, 0x2A, 0x3A, 0x55, 0x58, 0x13, 0x24, 0x21, 0x07, 0x5A, 0x3D, 0x69,
	0x1A, 0x0A, 0x09, 0x1A, 0x21, 0x3B, 0x35, 0x59, 0x09, 0x3A, 0x1F, 0x14,
	0x17, 0x31, 0x7A, 0x1C, 0x29, 0x05, 0x2C, 0x11, 0x3C, 0x51, 0x22, 0x3B,
	0x71, 0x1E, 0x28, 0x2C, 0x3B, 0x1A, 0x1F, 0x17, 0x18, 0x5E, 0x6D, 0x07,
	0x51, 0x38, 0x07, 0x69, 0x1A, 0x07, 0x26, 0x20, 0x7A, 0x04, 0x4E, 0x14,
	0x5D, 0x6D, 0x5D, 0x08, 0x59, 0x00, 0x6D, 0x58, 0x58, 0x34, 0x31, 0x75,
	0x35, 0x50, 0x58, 0x52, 0x2E, 0x1B, 0x26, 0x34, 0x0F, 0x72, 0x0D, 0x53,
	0x2B, 0x2F, 0x37, 0x08, 0x09, 0x3E, 0x1C, 0x26, 0x54, 0x59, 0x21, 0x52,
	0x24, 0x2E, 0x50, 0x57, 0x5B, 0x26, 0x09, 0x54, 0x21, 0x06, 0x20, 0x24,
	0x56, 0x2B, 0x19, 0x30, 0x28, 0x2C, 0x17, 0x19, 0x72, 0x0E, 0x53, 0x3C,
	0x52, 0x7B, 0x55, 0x04, 0x56, 0x13, 0x05, 0x1D, 0x3B, 0x0B, 0x24, 0x28,
	0x23, 0x33, 0x0A, 0x58, 0x05, 0x5E, 0x0A, 0x2C, 0x31, 0x28, 0x14, 0x16,
	0x5E, 0x24, 0x15, 0x01, 0x2D, 0x19, 0x5F, 0x01, 0x3B, 0x09, 0x2F, 0x1C,
	0x20, 0x24, 0x4E, 0x45, 0x3C, 0x30, 0x36, 0x52, 0x5C, 0x11, 0x15, 0x1C,
	0x24, 0x37, 0x3B, 0x35, 0x5C, 0x27, 0x1F, 0x05, 0x08, 0x0D, 0x58, 0x24,
	0x0D, 0x13, 0x19, 0x05, 0x06, 0x3C, 0x72, 0x1E, 0x18, 0x2F, 0x1F, 0x72,
	0x28, 0x0C, 0x0C, 0x05, 0x03, 0x01, 0x0B, 0x2C, 0x32, 0x31, 0x2B, 0x4A,
	0x14, 0x23, 0x29, 0x34, 0x26, 0x2D, 0x1A, 0x20, 0x0A, 0x0F, 0x5F, 0x12,
	0x72, 0x36, 0x30, 0x28, 0x24, 0x69, 0x01, 0x54, 0x2B, 0x31, 0x6D, 0x00,
	0x03, 0x20, 0x1C, 0x16, 0x14, 0x0E, 0x20, 0x28, 0x13, 0x1A, 0x0C, 0x00,
	0x5E, 0x12, 0x06, 0x3B, 0x0C, 0x12, 0x32, 0x29, 0x03, 0x3A, 0x1D, 0x04,
	0x3F, 0x2B, 0x03, 0x32, 0x1B, 0x0F, 0x00, 0x2A, 0x5B, 0x3B, 0x5C, 0x1B,
	0x06, 0x1F, 0x12, 0x29, 0x0D, 0x28, 0x12, 0x0E, 0x22, 0x4A, 0x00, 0x05,
	0x06, 0x3B, 0x28, 0x5D, 0x2D, 0x14, 0x02, 0x59, 0x38, 0x26, 0x0C, 0x23,
	0x39, 0x28, 0x33, 0x74, 0x3F, 0x2B, 0x27, 0x44, 0x26, 0x0F, 0x0E, 0x1A,
	0x5B, 0x07, 0x24, 0x36, 0x08, 0x2C, 0x77, 0x0B, 0x56, 0x1A, 0x3B, 0x24,
	0x5C, 0x17, 0x1D, 0x58, 0x2E, 0x24, 0x0E, 0x5D, 0x5A, 0x20, 0x23, 0x56,
	0x5B, 0x2A, 0x06, 0x5A, 0x04, 0x38, 0x33, 0x34, 0x23, 0x1B, 0x29, 0x0C,
	0x2C, 0x02, 0x4A, 0x0A, 0x3C, 0x0F, 0x54, 0x4E, 0x26, 0x1C, 0x36, 0x36,
	0x38, 0x24, 0x33, 0x0E, 0x1A, 0x27, 0x2B, 0x23, 0x2D, 0x35, 0x57, 0x02,
	0x44, 0x09, 0x5F, 0x2C, 0x28, 0x1C, 0x2A, 0x5E, 0x37, 0x17, 0x29, 0x70,
	0x00, 0x56, 0x3D, 0x0C, 0x2C, 0x15, 0x2C, 0x5D, 0x53, 0x71, 0x3B, 0x24,
	0x57, 0x3C, 0x74, 0x2D, 0x00, 0x23, 0x27, 0x3B, 0x0E, 0x2D, 0x5D, 0x0A,
	0x17, 0x3D, 0x2F, 0x23, 0x3B, 0x0F, 0x54, 0x4E, 0x27, 0x5D, 0x70, 0x43,
	0x17, 0x0F, 0x3F, 0x7A, 0x28, 0x59, 0x1A, 0x06, 0x25, 0x20, 0x16, 0x01,
	0x44, 0x6D, 0x09, 0x31, 0x5E, 0x09, 0x12, 0x5E, 0x57, 0x05, 0x5F, 0x11,
	0x5D, 0x51, 0x04, 0x26, 0x20, 0x43, 0x11, 0x1B, 0x53, 0x21, 0x02, 0x2B,
	0x1B, 0x2C, 0x2F, 0x34, 0x29, 0x41, 0x24, 0x20, 0x5B, 0x0A, 0x1F, 0x2F,
	0x14, 0x21, 0x0E, 0x5D, 0x3A, 0x1A, 0x01, 0x06, 0x38, 0x2D, 0x16, 0x20,
	0x54, 0x22, 0x40, 0x70, 0x09, 0x11, 0x1D, 0x00, 0x0D, 0x00, 0x17, 0x38,
	0x2D, 0x71, 0x2F, 0x37, 0x5F, 0x27, 0x7A, 0x25, 0x4A, 0x21, 0x39, 0x0D,
	0x15, 0x2E, 0x05, 0x07, 0x37, 0x2B, 0x37, 0x39, 0x0D, 0x23, 0x38, 0x12,
	0x3E, 0x28, 0x28, 0x00, 0x02, 0x21, 0x09, 0x0D, 0x1A, 0x34, 0x06, 0x53,
	0x1B, 0x58, 0x15, 0x58, 0x5F, 0x3A, 0x05, 0x59, 0x00, 0x1C, 0x70, 0x08,
	0x19, 0x36, 0x5F, 0x0D, 0x14, 0x36, 0x28, 0x0E, 0x6D, 0x20, 0x3B, 0x2F,
	0x1C, 0x76, 0x54, 0x18, 0x1F, 0x2F, 0x7A, 0x0E, 0x02, 0x5F, 0x31, 0x2A,
	0x2E, 0x11, 0x16, 0x23, 0x2F, 0x5D, 0x37, 0x08, 0x00, 0x21, 0x34, 0x02,
	0x5C, 0x20, 0x34, 0x04, 0x22, 0x45, 0x22, 0x2C, 0x3C, 0x34, 0x1F, 0x11,
	0x72, 0x2B, 0x34, 0x36, 0x1E, 0x74, 0x38, 0x32, 0x57, 0x24, 0x3A, 0x1A,
	0x23, 0x23, 0x25, 0x08, 0x0F, 0x07, 0x2B, 0x0C, 0x26, 0x2D, 0x54, 0x02,
	0x3A, 0x18, 0x2B, 0x10, 0x23, 0x2E, 0x31, 0x23, 0x51, 0x3B, 0x1A, 0x0A,
	0x2D, 0x06, 0x45, 0x1B, 0x34, 0x5E, 0x0E, 0x5F, 0x2C, 0x01, 0x03, 0x53,
	0x3B, 0x5E, 0x2A, 0x2E, 0x13, 0x26, 0x5F, 0x1B, 0x34, 0x00, 0x36, 0x5D,
	0x71, 0x15, 0x2D, 0x59, 0x2E, 0x30, 0x14, 0x06, 0x05, 0x29, 0x71, 0x02,
	0x31, 0x1F, 0x5C, 0x27, 0x22, 0x33, 0x1F, 0x5E, 0x6D, 0x1E, 0x09, 0x2A,
	0x58, 0x33, 0x20, 0x04, 0x2D, 0x32, 0x69, 0x0B, 0x11, 0x56, 0x18, 0x36,
	0x5C, 0x13, 0x3E, 0x02, 0x0A, 0x43, 0x23, 0x58, 0x06, 0x75, 0x25, 0x51,
	0x0A, 0x25, 0x14, 0x15, 0x2C, 0x3C, 0x19, 0x3B, 0x58, 0x0A, 0x5A, 0x2D,
	0x0D, 0x05, 0x50, 0x28, 0x23, 0x38, 0x21, 0x51, 0x5E, 0x3D, 0x00, 0x21,
	0x0D, 0x5E, 0x22, 0x05, 0x2B, 0x0F, 0x2D, 0x05, 0x04, 0x29, 0x59, 0x24,
	0x5D, 0x15, 0x0E, 0x12, 0x0B, 0x23, 0x33, 0x05, 0x0D, 0x2C, 0x32, 0x14,
	0x38, 0x04, 0x1E, 0x28, 0x26, 0x06, 0x28, 0x27, 0x2D, 0x7A, 0x20, 0x37,
	0x5C, 0x12, 0x0D, 0x5C, 0x16, 0x1C, 0x20, 0x23, 0x34, 0x0E, 0x1E, 0x31,
	0x35, 0x25, 0x0F, 0x1C, 0x20, 0x03, 0x59, 0x2F, 0x38, 0x25, 0x01, 0x3C,
	0x08, 0x23, 0x08, 0x31, 0x27, 0x33, 0x5A, 0x11, 0x27, 0x1D, 0x2C, 0x1F,
	0x01, 0x26, 0x02, 0x0D, 0x16, 0x22, 0x3A, 0x14, 0x0C, 0x07, 0x2C, 0x0F,
	0x0E, 0x22, 0x07, 0x33, 0x74, 0x0F, 0x04, 0x3C, 0x00, 0x34, 0x3D, 0x31,
	0x1D, 0x09, 0x05, 0x29, 0x4A, 0x3F, 0x07, 0x10, 0x0E, 0x56, 0x23, 0x1C,
	0x0B, 0x43, 0x55, 0x0F, 0x00, 0x30, 0x1D, 0x2D, 0x5D, 0x09, 0x2F, 0x00,
	0x59, 0x22, 0x0D, 0x24, 0x59, 0x50, 0x17, 0x25, 0x35, 0x29, 0x55, 0x38,
	0x5A, 0x0E, 0x26, 0x0D, 0x57, 0x03, 0x21, 0x03, 0x30, 0x23, 0x1C, 0x23,
	0x20, 0x2C, 0x00, 0x3F, 0x1B, 0x09, 0x03, 0x14, 0x38, 0x75, 0x23, 0x38,
	0x0A, 0x09, 0x36, 0x2A, 0x04, 0x56, 0x32, 0x1B, 0x54, 0x1B, 0x1D, 0x2D,
	0x04, 0x3A, 0x2F, 0x00, 0x1C, 0x1A, 0x02, 0x34, 0x5A, 0x03, 0x38, 0x20,
	0x20, 0x3D, 0x3B, 0x69, 0x06, 0x09, 0x01, 0x3B, 0x34, 0x43, 0x2B, 0x03,
	0x3C, 0x31, 0x08, 0x17, 0x34, 0x04, 0x15, 0x29, 0x4A, 0x21, 0x1E, 0x2D,
	0x09, 0x31, 0x2C, 0x5D, 0x34, 0x3A, 0x57, 0x17, 0x2D, 0x70, 0x06, 0x23,
	0x00, 0x11, 0x77, 0x08, 0x16, 0x16, 0x5F, 0x70, 0x39, 0x24, 0x28, 0x2D,
	0x74, 0x55, 0x50, 0x37, 0x26, 0x32, 0x36, 0x3B, 0x41, 0x59, 0x1B, 0x15,
	0x1B, 0x16, 0x2C, 0x36, 0x2B, 0x18, 0x06, 0x44, 0x74, 0x21, 0x55, 0x0C,
	0x09, 0x73, 0x3E, 0x0B, 0x08, 0x1E, 0x15, 0x3D, 0x14, 0x09, 0x2D, 0x14,
	0x22, 0x03, 0x3F, 0x3B, 0x09, 0x03, 0x52, 0x38, 0x0A, 0x35, 0x19, 0x13,
	0x3D, 0x2A, 0x0D, 0x5D, 0x4E, 0x0A, 0x59, 0x77, 0x18, 0x11, 0x3E, 0x38,
	0x23, 0x5F, 0x32, 0x06, 0x27, 0x21, 0x36, 0x20, 0x27, 0x1D, 0x15, 0x59,
	0x03, 0x00, 0x27, 0x7B, 0x0D, 0x26, 0x20, 0x0A, 0x06, 0x14, 0x10, 0x01,
	0x5A, 0x37, 0x22, 0x56, 0x09, 0x1D, 0x07, 0x28, 0x31, 0x2A, 0x01, 0x3A,
	0x35, 0x4E, 0x58, 0x31, 0x28, 0x06, 0x17, 0x01, 0x1F, 0x23, 0x58, 0x0A,
	0x57, 0x0A, 0x28, 0x38, 0x2D, 0x03, 0x31, 0x71, 0x2A, 0x09, 0x56, 0x38,
	0x70, 0x29, 0x27, 0x04, 0x1D, 0x09, 0x2E, 0x58, 0x18, 0x44, 0x2D, 0x08,
	0x35, 0x25, 0x04, 0x74, 0x5E, 0x4A, 0x08, 0x3D, 0x09, 0x28, 0x02, 0x24,
	0x5D, 0x03, 0x06, 0x09, 0x29, 0x5A, 0x3A, 0x2B, 0x2D, 0x27, 0x23, 0x18,
	0x5C, 0x52, 0x2B, 0x52, 0x1A, 0x04, 0x20, 0x0A, 0x2A, 0x33, 0x3E, 0x04,
	0x3A, 0x29, 0x35, 0x29, 0x51, 0x17, 0x19, 0x73, 0x54, 0x55, 0x18, 0x02,
	0x38, 0x20, 0x35, 0x00, 0x22, 0x2D, 0x24, 0x05, 0x37, 0x22, 0x30, 0x2B,
	0x31, 0x14, 0x0C, 0x21, 0x1D, 0x0E, 0x16, 0x19, 0x2A, 0x04, 0x32, 0x14,
	0x5D, 0x11, 0x00, 0x19, 0x2A, 0x03, 0x23, 0x1E, 0x2F, 0x01, 0x2D, 0x73,
	0x20, 0x28, 0x16, 0x5A, 0x1A, 0x0B, 0x05, 0x38, 0x2D, 0x73, 0x19, 0x07,
	0x1F, 0x1F, 0x10, 0x0D, 0x11, 0x38, 0x0E, 0x25, 0x5F, 0x0E, 0x04, 0x5D,
	0x72, 0x01, 0x0E, 0x22, 0x24, 0x75, 0x5A, 0x25, 0x41, 0x52, 0x13, 0x16,
	0x33, 0x5D, 0x2A, 0x0B, 0x23, 0x51, 0x5A, 0x26, 0x10, 0x07, 0x0F, 0x2F,
	0x5E, 0x00, 0x26, 0x54, 0x04, 0x21, 0x04, 0x25, 0x59, 0x05, 0x12, 0x38,
	0x09, 0x06, 0x5D, 0x07, 0x20, 0x28, 0x2F, 0x38, 0x32, 0x2D, 0x1B, 0x31,
	0x2B, 0x2C, 0x0C, 0x1E, 0x32, 0x0A, 0x5F, 0x15, 0x1F, 0x58, 0x58, 0x00,
	0x03, 0x1E, 0x37, 0x0D, 0x1A, 0x10, 0x2E, 0x0F, 0x58, 0x02, 0x16, 0x2B,
	0x35, 0x09, 0x13, 0x25, 0x04, 0x2B, 0x1E, 0x2E, 0x00, 0x01, 0x2D, 0x0D,
	0x26, 0x72, 0x16, 0x2C, 0x03, 0x18, 0x76, 0x35, 0x57, 0x20, 0x32, 0x29,
	0x43, 0x35, 0x16, 0x1F, 0x11, 0x39, 0x14, 0x14, 0x5B, 0x7A, 0x3E, 0x14,
	0x2F, 0x13, 0x32, 0x1A, 0x11, 0x2F, 0x0C, 0x77, 0x19, 0x59, 0x21, 0x26,
	0x28, 0x54, 0x2B, 0x06, 0x22, 0x74, 0x19, 0x14, 0x2A, 0x31, 0x10, 0x34,
	0x32, 0x28, 0x22, 0x34, 0x16, 0x06, 0x3D, 0x52, 0x0D, 0x29, 0x25, 0x5E,
	0x2D, 0x30, 0x5E, 0x2A, 0x1D, 0x3D, 0x27, 0x21, 0x10, 0x57, 0x3F, 0x3B,
	0x39, 0x34, 0x25, 0x08, 0x7B, 0x14, 0x2B, 0x5A, 0x5C, 0x2B, 0x5D, 0x58,
	0x0D, 0x59, 0x2E, 0x1F, 0x0F, 0x20, 0x18, 0x11, 0x23, 0x31, 0x5C, 0x1F,
	0x2A, 0x25, 0x1B, 0x0B, 0x29, 0x75, 0x00, 0x02, 0x0F, 0x1F, 0x0A, 0x1D,
	0x09, 0x3E, 0x5C, 0x73, 0x07, 0x04, 0x3E, 0x1A, 0x69, 0x2A, 0x29, 0x3B,
	0x53, 0x36, 0x34, 0x50, 0x2F, 0x18, 0x0F, 0x3B, 0x09, 0x1F, 0x1F, 0x70,
	0x07, 0x55, 0x56, 0x26, 0x72, 0x58, 0x50, 0x5D, 0x5D, 0x30, 0x5C, 0x02,
	0x29, 0x1E, 0x73, 0x39, 0x30, 0x1F, 0x3E, 0x2C, 0x22, 0x27, 0x08, 0x20,
	0x03, 0x05, 0x29, 0x0B, 0x27, 0x0D, 0x03, 0x25, 0x06, 0x5A, 0x07, 0x5C,
	0x13, 0x07, 0x26, 0x74, 0x2B, 0x12, 0x3F, 0x04, 0x2D, 0x5D, 0x30, 0x0D,
	0x00, 0x05, 0x2D, 0x53, 0x17, 0x1A, 0x25, 0x2A, 0x4A, 0x14, 0x1F, 0x01,
	0x05, 0x58, 0x58, 0x0C, 0x29, 0x14, 0x2C, 0x0F, 0x2D, 0x2A, 0x5C, 0x52,
	0x5A, 0x2F, 0x36, 0x5B, 0x07, 0x17, 0x25, 0x28, 0x25, 0x54, 0x14, 0x2E,
	0x31, 0x03, 0x52, 0x36, 0x5D, 0x24, 0x28, 0x05, 0x3D, 0x3C, 0x3B, 0x3A,
	0x18, 0x34, 0x3F, 0x37, 0x3D, 0x13, 0x16, 0x26, 0x38, 0x59, 0x0D, 0x0C,
	0x19, 0x0A, 0x5B, 0x39, 0x2D, 0x0E, 0x0B, 0x0E, 0x55, 0x04, 0x21, 0x0A,
	0x2A, 0x59, 0x0A, 0x21, 0x06, 0x04, 0x33, 0x04, 0x3A, 0x0F, 0x38, 0x20,
	0x18, 0x18, 0x7A, 0x21, 0x20, 0x06, 0x0E, 0x1A, 0x59, 0x39, 0x1F, 0x00,
	0x2A, 0x27, 0x2F, 0x1B, 0x11, 0x20, 0x03, 0x19, 0x26, 0x3D, 0x20, 0x00,
	0x03, 0x1B, 0x19, 0x1A, 0x16, 0x2C, 0x2C, 0x25, 0x0C, 0x35, 0x54, 0x05,
	0x3A, 0x2B, 0x3A, 0x08, 0x5E, 0x3B, 0x31, 0x5C, 0x14, 0x41, 0x1C, 0x04,
	0x3B, 0x0B, 0x57, 0x53, 0x20, 0x1E, 0x0C, 0x17, 0x33, 0x32, 0x0F, 0x13,
	0x19, 0x5A, 0x2B, 0x2A, 0x52, 0x19, 0x5F, 0x14, 0x34, 0x0C, 0x22, 0x1B,
	0x2C, 0x29, 0x00, 0x00, 0x02, 0x70, 0x26, 0x33, 0x0F, 0x59, 0x0D, 0x3A,
	0x34, 0x00, 0x0D, 0x37, 0x22, 0x25, 0x0C, 0x04, 0x23, 0x3A, 0x1B, 0x27,
	0x5B, 0x2B, 0x05, 0x23, 0x20, 0x24, 0x74, 0x16, 0x55, 0x2C, 0x00, 0x29,
	0x2A, 0x31, 0x41, 0x04, 0x76, 0x5A, 0x05, 0x17, 0x28, 0x35, 0x58, 0x2E,
	0x56, 0x3C, 0x17, 0x3D, 0x3B, 0x45, 0x13, 0x09, 0x05, 0x50, 0x21, 0x23,
	0x7A, 0x25, 0x0E, 0x1A, 0x0D, 0x06, 0x1C, 0x59, 0x07, 0x25, 0x70, 0x19,
	0x3B, 0x0D, 0x25, 0x26, 0x06, 0x2C, 0x03, 0x38, 0x30, 0x27, 0x26, 0x21,
	0x32, 0x11, 0x08, 0x1B, 0x1A, 0x59, 0x20, 0x3B, 0x03, 0x22, 0x3A, 0x77,
	0x3B, 0x31, 0x2F, 0x07, 0x1B, 0x54, 0x0A, 0x07, 0x40, 0x0A, 0x34, 0x13,
	0x3C, 0x40, 0x12, 0x0F, 0x59, 0x03, 0x04, 0x74, 0x43, 0x51, 0x0F, 0x09,
	0x2B, 0x07, 0x2B, 0x07, 0x53, 0x35, 0x29, 0x39, 0x3A, 0x04, 0x75, 0x14,
	0x0D, 0x2A, 0x59, 0x15, 0x3A, 0x3B, 0x18, 0x0E, 0x0B, 0x1E, 0x2C, 0x28,
	0x1D, 0x18, 0x47, 0x16, 0x23, 0x58, 0x75, 0x1E, 0x18, 0x2B, 0x00, 0x32,
	0x5E, 0x55, 0x00, 0x38, 0x12, 0x36, 0x3B, 0x07, 0x29, 0x38, 0x0E, 0x0E,
	0x5F, 0x2C, 0x20, 0x3B, 0x07, 0x1B, 0x1F, 0x3B, 0x5C, 0x52, 0x3D, 0x40,
	0x2B, 0x20, 0x20, 0x39, 0x33, 0x29, 0x5C, 0x26, 0x09, 0x29, 0x08, 0x59,
	0x0D, 0x5F, 0x27, 0x15, 0x5A, 0x37, 0x17, 0x11, 0x25, 0x3F, 0x0E, 0x0C,
	0x25, 0x3A, 0x07, 0x59, 0x0F, 0x28, 0x72, 0x5F, 0x36, 0x59, 0x38, 0x37,
	0x1C, 0x52, 0x0C, 0x2A, 0x07, 0x58, 0x57, 0x23, 0x0C, 0x2C, 0x2B, 0x03,
	0x03, 0x1D, 0x08, 0x54, 0x2F, 0x26, 0x04, 0x11, 0x2B, 0x58, 0x0B, 0x28,
	0x2A, 0x36, 0x13, 0x41, 0x03, 0x14, 0x24, 0x0F, 0x09, 0x33, 0x0A, 0x5F,
	0x16, 0x17, 0x25, 0x2F, 0x02, 0x52, 0x39, 0x06, 0x7B, 0x0D, 0x16, 0x14,
	0x01, 0x10, 0x54, 0x09, 0x16, 0x3B, 0x31, 0x23, 0x0D, 0x0F, 0x00, 0x2B,
	0x3A, 0x0E, 0x3D, 0x0A, 0x00, 0x2E, 0x24, 0x41, 0x04, 0x04, 0x5D, 0x38,
	0x0A, 0x5A, 0x36, 0x1D, 0x3B, 0x09, 0x5A, 0x38, 0x23, 0x39, 0x3C, 0x5C,
	0x2B, 0x5D, 0x00, 0x07, 0x40, 0x38, 0x3C, 0x2A, 0x1B, 0x3B, 0x72, 0x02,
	0x33, 0x56, 0x24, 0x7B, 0x55, 0x18, 0x3D, 0x26, 0x2A, 0x07, 0x34, 0x0F,
	0x01, 0x1B, 0x0D, 0x57, 0x09, 0x26, 0x31, 0x15, 0x00, 0x2B, 0x0E, 0x74,
	0x35, 0x52, 0x34, 0x1B, 0x2F, 0x06, 0x11, 0x59, 0x29, 0x0B, 0x5C, 0x56,
	0x05, 0x40, 0x2D, 0x43, 0x0B, 0x45, 0x3D, 0x6D, 0x58, 0x11, 0x41, 0x0C,
	0x0F, 0x39, 0x27, 0x2F, 0x13, 0x07, 0x39, 0x29, 0x0F, 0x12, 0x07, 0x1F,
	0x09, 0x2B, 0x53, 0x1B, 0x25, 0x25, 0x0D, 0x59, 0x31, 0x23, 0x59, 0x3B,
	0x33, 0x06, 0x2E, 0x20, 0x36, 0x07, 0x10, 0x14, 0x59, 0x07, 0x21, 0x18,
	0x5E, 0x52, 0x29, 0x0A, 0x24, 0x38, 0x07, 0x06, 0x09, 0x29, 0x1E, 0x2B,
	0x59, 0x31, 0x69, 0x35, 0x07, 0x57, 0x39, 0x2D, 0x27, 0x24, 0x2A, 0x03,
	0x6D, 0x06, 0x26, 0x01, 0x0D, 0x03, 0x5F, 0x00, 0x29, 0x3E, 0x12, 0x43,
	0x51, 0x0D, 0x53, 0x01, 0x09, 0x38, 0x1D, 0x27, 0x36, 0x14, 0x51, 0x16,
	0x2A, 0x09, 0x55, 0x56, 0x20, 0x08, 0x10, 0x5D, 0x53, 0x1A, 0x0C, 0x36,
	0x5E, 0x38, 0x59, 0x04, 0x32, 0x5D, 0x2B, 0x24, 0x39, 0x0E, 0x01, 0x33,
	0x3C, 0x04, 0x3A, 0x43, 0x0E, 0x14, 0x38, 0x13, 0x54, 0x37, 0x22, 0x04,
	0x31, 0x00, 0x0A, 0x28, 0x53, 0x2C, 0x5A, 0x39, 0x1C, 0x24, 0x23, 0x5D,
	0x55, 0x5A, 0x05, 0x0A, 0x09, 0x29, 0x1C, 0x13, 0x73, 0x2B, 0x53, 0x16,
	0x2A, 0x21, 0x03, 0x22, 0x2D, 0x3F, 0x13, 0x0E, 0x07, 0x5E, 0x31, 0x30,
	0x18, 0x53, 0x5A, 0x04, 0x25, 0x24, 0x56, 0x5F, 0x2F, 0x1A, 0x03, 0x14,
	0x19, 0x32, 0x1A, 0x2A, 0x08, 0x5E, 0x2D, 0x2C, 0x07, 0x0C, 0x22, 0x05,
	0x74, 0x59, 0x13, 0x27, 0x5D, 0x07, 0x1C, 0x32, 0x23, 0x19, 0x24, 0x09,
	0x2B, 0x06, 0x01, 0x17, 0x1A, 0x52, 0x5B, 0x01, 0x0F, 0x22, 0x30, 0x19,
	0x44, 0x24, 0x34, 0x36, 0x45, 0x06, 0x0B, 0x35, 0x59, 0x0B, 0x20, 0x2C,
	0x36, 0x37, 0x56, 0x1C, 0x3A, 0x5F, 0x34, 0x01, 0x01, 0x3A, 0x5E, 0x15,
	0x5A, 0x5C, 0x74, 0x2B, 0x55, 0x37, 0x40, 0x70, 0x36, 0x59, 0x21, 0x00,
	0x0D, 0x38, 0x53, 0x0F, 0x3C, 0x7B, 0x16, 0x30, 0x02, 0x53, 0x35, 0x15,
	0x55, 0x1D, 0x2C, 0x34, 0x5C, 0x33, 0x28, 0x0F, 0x29, 0x04, 0x2D, 0x21,
	0x58, 0x0C, 0x07, 0x12, 0x34, 0x12, 0x27, 0x05, 0x2E, 0x08, 0x18, 0x75,
	0x1D, 0x34, 0x00, 0x00, 0x30, 0x08, 0x26, 0x0D, 0x0D, 0x7A, 0x20, 0x0B,
	0x1F, 0x38, 0x73, 0x2B, 0x12, 0x39, 0x1A, 0x20, 0x25, 0x32, 0x26, 0x44,
	0x74, 0x25, 0x04, 0x59, 0x33, 0x2E, 0x55, 0x52, 0x19, 0x22, 0x30, 0x2E,
	0x51, 0x36, 0x5B, 0x16, 0x43, 0x2A, 0x41, 0x2A, 0x3B, 0x1F, 0x24, 0x0A,
	0x05, 0x2F, 0x04, 0x2E, 0x57, 0x38, 0x07, 0x06, 0x25, 0x22, 0x52, 0x20,
	0x26, 0x36, 0x56, 0x58, 0x28, 0x2D, 0x53, 0x1C, 0x2F, 0x15, 0x1B, 0x24,
	0x22, 0x5C, 0x20, 0x0B, 0x0C, 0x2B, 0x52, 0x71, 0x34, 0x0E, 0x37, 0x03,
	0x06, 0x0A, 0x06, 0x58, 0x5E, 0x0F, 0x47, 0x22, 0x3B, 0x26, 0x12, 0x34,
	0x29, 0x09, 0x18, 0x20, 0x27, 0x0B, 0x5C, 0x3C, 0x05, 0x2D, 0x31, 0x5E,
	0x22, 0x32, 0x15, 0x15, 0x19, 0x59, 0x28, 0x23, 0x04, 0x23, 0x01, 0x0C,
	0x5D, 0x2E, 0x04, 0x2D, 0x72, 0x27, 0x06, 0x1C, 0x20, 0x6D, 0x2B, 0x35,
	0x5F, 0x40, 0x2F, 0x5D, 0x2C, 0x06, 0x1D, 0x34, 0x5E, 0x1B, 0x5F, 0x0C,
	0x1B, 0x22, 0x56, 0x02, 0x04, 0x03, 0x0B, 0x2E, 0x39, 0x3D, 0x1A, 0x22,
	0x15, 0x2A, 0x03, 0x04, 0x3E, 0x18, 0x00, 0x27, 0x72, 0x3C, 0x11, 0x38,
	0x02, 0x69, 0x0D, 0x51, 0x0F, 0x3E, 0x18, 0x28, 0x54, 0x17, 0x01, 0x3B,
	0x09, 0x52, 0x1F, 0x28, 0x11, 0x26, 0x27, 0x21, 0x3B, 0x18, 0x22, 0x28,
	0x24, 0x53, 0x2C, 0x34, 0x32, 0x18, 0x27, 0x11, 0x22, 0x23, 0x3C, 0x2F,
	0x15, 0x25, 0x2F, 0x23, 0x2F, 0x05, 0x29, 0x05, 0x57, 0x13, 0x7B, 0x5D,
	0x35, 0x20, 0x3F, 0x0A, 0x5C, 0x34, 0x2B, 0x18, 0x17, 0x15, 0x2F, 0x19,
	0x1A, 0x04, 0x23, 0x0C, 0x18, 0x1D, 0x21, 0x1E, 0x18, 0x23, 0x05, 0x16,
	0x36, 0x54, 0x06, 0x3E, 0x29, 0x00, 0x20, 0x3F, 0x59, 0x14, 0x2A, 0x31,
	0x27, 0x27, 0x7A, 0x0E, 0x04, 0x2D, 0x09, 0x26, 0x58, 0x0E, 0x37, 0x1A,
	0x01, 0x36, 0x57, 0x16, 0x1A, 0x07, 0x23, 0x4E, 0x19, 0x0E, 0x74, 0x2F,
	0x26, 0x3B, 0x25, 0x71, 0x16, 0x0D, 0x3D, 0x33, 0x73, 0x0D, 0x07, 0x25,
	0x19, 0x77, 0x1B, 0x0F, 0x22, 0x01, 0x2D, 0x2A, 0x4E, 0x19, 0x3B, 0x38,
	0x14, 0x2F, 0x57, 0x2E, 0x09, 0x1F, 0x59, 0x0D, 0x25, 0x1B, 0x5F, 0x10,
	0x22, 0x09, 0x37, 0x2E, 0x12, 0x00, 0x5D, 0x27, 0x04, 0x0A, 0x5F, 0x12,
	0x75, 0x38, 0x19, 0x16, 0x5A, 0x7B, 0x25, 0x51, 0x59, 0x08, 0x74, 0x03,
	0x07, 0x06, 0x53, 0x24, 0x0F, 0x2B, 0x45, 0x5C, 0x77, 0x2E, 0x30, 0x17,
	0x5F, 0x04, 0x3B, 0x29, 0x56, 0x27, 0x00, 0x27, 0x23, 0x2D, 0x5A, 0x09,
	0x3D, 0x00, 0x45, 0x3D, 0x25, 0x5E, 0x13, 0x2A, 0x0E, 0x13, 0x26, 0x04,
	0x5D, 0x44, 0x0C, 0x16, 0x51, 0x22, 0x32, 0x74, 0x43, 0x19, 0x59, 0x27,
	0x0E, 0x15, 0x51, 0x0D, 0x1E, 0x77, 0x3A, 0x2B, 0x04, 0x52, 0x76, 0x05,
	0x26, 0x20, 0x5E, 0x2E, 0x06, 0x08, 0x1E, 0x1E, 0x74, 0x0F, 0x33, 0x5C,
	0x59, 0x2A, 0x20, 0x1B, 0x22, 0x5D, 0x33, 0x5A, 0x51, 0x3C, 0x05, 0x77,
	0x0A, 0x13, 0x0F, 0x53, 0x0F, 0x43, 0x34, 0x56, 0x31, 0x09, 0x09, 0x15,
	0x22, 0x07, 0x3B, 0x02, 0x31, 0x18, 0x21, 0x76, 0x04, 0x56, 0x34, 0x00,
	0x76, 0x23, 0x50, 0x37, 0x5D, 0x07, 0x47, 0x08, 0x08, 0x05, 0x24, 0x26,
	0x06, 0x3E, 0x3B, 0x23, 0x25, 0x55, 0x0C, 0x2E, 0x0D, 0x08, 0x23, 0x39,
	0x32, 0x33, 0x28, 0x1B, 0x5C, 0x1D, 0x1B, 0x3F, 0x4E, 0x0C, 0x12, 0x70,
	0x1C, 0x51, 0x3F, 0x44, 0x30, 0x5D, 0x50, 0x0D, 0x04, 0x32, 0x43, 0x39,
	0x22, 0x06, 0x17, 0x3C, 0x2D, 0x45, 0x39, 0x15, 0x1F, 0x20, 0x0D, 0x32,
	0x14, 0x18, 0x0B, 0x2A, 0x03, 0x36, 0x14, 0x00, 0x57, 0x1D, 0x00, 0x3B,
	0x03, 0x06, 0x5A, 0x75, 0x5E, 0x2B, 0x19, 0x09, 0x25, 0x2D, 0x07, 0x5B,
	0x3A, 0x72, 0x02, 0x04, 0x3D, 0x09, 0x21, 0x0A, 0x32, 0x2B, 0x19, 0x0D,
	0x2A, 0x3B, 0x1A, 0x13, 0x0B, 0x5F, 0x2B, 0x57, 0x19, 0x2F, 0x5C, 0x57,
	0x1C, 0x04, 0x34, 0x02, 0x57, 0x26, 0x20, 0x08, 0x1F, 0x14, 0x59, 0x59,
	0x16, 0x5A, 0x51, 0x01, 0x1B, 0x33, 0x1A, 0x00, 0x5F, 0x2D, 0x34, 0x1C,
	0x4A, 0x22, 0x00, 0x7B, 0x5D, 0x14, 0x5E, 0x00, 0x12, 0x25, 0x56, 0x1D,
	0x3E, 0x1B, 0x09, 0x14, 0x24, 0x0F, 0x05, 0x5C, 0x0A, 0x27, 0x5B, 0x15,
	0x24, 0x0B, 0x28, 0x19, 0x12, 0x25, 0x56, 0x38, 0x5B, 0x18, 0x16, 0x0D,
	0x1F, 0x1B, 0x0A, 0x5D, 0x37, 0x0A, 0x00, 0x17, 0x5F, 0x36, 0x5C, 0x2E,
	0x69, 0x1A, 0x0A, 0x3A, 0x3D, 0x30, 0x15, 0x32, 0x03, 0x3A, 0x16, 0x0A,
	0x34, 0x01, 0x5A, 0x33, 0x24, 0x50, 0x1A, 0x5C, 0x3A, 0x43, 0x27, 0x58,
	0x0E, 0x2D, 0x1B, 0x11, 0x22, 0x40, 0x38, 0x29, 0x34, 0x0F, 0x3C, 0x06,
	0x1E, 0x0E, 0x26, 0x40, 0x0D, 0x39, 0x35, 0x5D, 0x18, 0x77, 0x0A, 0x37,
	0x09, 0x0E, 0x15, 0x5F, 0x32, 0x08, 0x5D, 0x32, 0x43, 0x59, 0x2B, 0x2E,
	0x7A, 0x08, 0x13, 0x0B, 0x5D, 0x05, 0x0F, 0x16, 0x1B, 0x31, 0x7A, 0x26,
	0x10, 0x34, 0x2C, 0x20, 0x08, 0x2A, 0x3A, 0x0E, 0x73, 0x0A, 0x20, 0x0A,
	0x03, 0x24, 0x0F, 0x29, 0x2F, 0x26, 0x14, 0x3B, 0x0E, 0x29, 0x2F, 0x75,
	0x2E, 0x56, 0x1A, 0x1C, 0x36, 0x3F, 0x36, 0x01, 0x2F, 0x31, 0x09, 0x22,
	0x24, 0x38, 0x17, 0x29, 0x11, 0x21, 0x31, 0x25, 0x1B, 0x39, 0x24, 0x28,
	0x00, 0x43, 0x36, 0x20, 0x2A, 0x0E, 0x0F, 0x18, 0x23, 0x3A, 0x0F, 0x27,
	0x26, 0x0D, 0x5B, 0x77, 0x2E, 0x29, 0x20, 0x04, 0x21, 0x1E, 0x38, 0x1A,
	0x20, 0x18, 0x23, 0x53, 0x5D, 0x12, 0x32, 0x3D, 0x0B, 0x19, 0x1E, 0x29,
	0x58, 0x07, 0x5F, 0x19, 0x10, 0x59, 0x0B, 0x02, 0x3F, 0x73, 0x29, 0x19,
	0x39, 0x0D, 0x74, 0x0F, 0x04, 0x09, 0x5E, 0x11, 0x18, 0x27, 0x20, 0x26,
	0x05, 0x2B, 0x18, 0x26, 0x00, 0x2F, 0x06, 0x26, 0x5F, 0x52, 0x24, 0x04,
	0x00, 0x5D, 0x07, 0x23, 0x01, 0x11, 0x06, 0x07, 0x0C, 0x58, 0x2C, 0x01,
	0x1D, 0x3A, 0x59, 0x06, 0x3D, 0x13, 0x0E, 0x1E, 0x54, 0x0A, 0x3B, 0x0F,
	0x39, 0x12, 0x1D, 0x5B, 0x34, 0x22, 0x13, 0x38, 0x04, 0x03, 0x5B, 0x39,
	0x2B, 0x5C, 0x12, 0x2E, 0x00, 0x14, 0x1B, 0x76, 0x2D, 0x22, 0x03, 0x40,
	0x7B, 0x36, 0x16, 0x3F, 0x38, 0x7A, 0x3F, 0x00, 0x05, 0x2E, 0x25, 0x21,
	0x12, 0x5F, 0x3A, 0x25, 0x2E, 0x20, 0x0D, 0x18, 0x72, 0x5A, 0x37, 0x27,
	0x2A, 0x23, 0x02, 0x3B, 0x39, 0x39, 0x25, 0x5A, 0x37, 0x23, 0x1B, 0x2E,
	0x07, 0x02, 0x14, 0x1A, 0x0D, 0x58, 0x05, 0x34, 0x5F, 0x2F, 0x22, 0x2B,
	0x0B, 0x5A, 0x76, 0x54, 0x57, 0x18, 0x09, 0x1B, 0x3E, 0x52, 0x2A, 0x09,
	0x69, 0x0B, 0x0E, 0x39, 0x06, 0x12, 0x21, 0x4E, 0x16, 0x0D, 0x05, 0x1A,
	0x25, 0x0F, 0x31, 0x0A, 0x19, 0x0E, 0x1D, 0x3E, 0x12, 0x15, 0x09, 0x03,
	0x38, 0x10, 0x36, 0x2C, 0x3B, 0x18, 0x38, 0x15, 0x53, 0x21, 0x2E, 0x1A,
	0x01, 0x0D, 0x3B, 0x1A, 0x2A, 0x18, 0x58, 0x3D, 0x26, 0x23, 0x19, 0x22,
	0x14, 0x01, 0x2A, 0x07, 0x4A, 0x39, 0x19, 0x32, 0x1C, 0x57, 0x25, 0x24,
	0x24, 0x01, 0x0E, 0x2D, 0x2F, 0x0B, 0x34, 0x38, 0x1B, 0x11, 0x00, 0x28,
	0x2E, 0x2B, 0x0A, 0x30, 0x3A, 0x4A, 0x05, 0x31, 0x0D, 0x0A, 0x35, 0x1C,
	0x44, 0x25, 0x16, 0x0A, 0x26, 0x3B, 0x29, 0x5D, 0x3B, 0x3D, 0x2F, 0x16,
	0x5D, 0x2B, 0x56, 0x29, 0x24, 0x2D, 0x58, 0x08, 0x26, 0x75, 0x23, 0x17,
	0x5A, 0x03, 0x24, 0x18, 0x19, 0x08, 0x2C, 0x34, 0x3A, 0x04, 0x06, 0x0D,
	0x72, 0x5D, 0x34, 0x07, 0x5B, 0x3A, 0x09, 0x2C, 0x5C, 0x26, 0x09, 0x15,
	0x37, 0x56, 0x25, 0x3B, 0x20, 0x34, 0x26, 0x1E, 0x24, 0x2F, 0x16, 0x41,
	0x1D, 0x2C, 0x22, 0x0A, 0x5B, 0x24, 0x69, 0x08, 0x2D, 0x2D, 0x25, 0x34,
	0x14, 0x0B, 0x25, 0x02, 0x24, 0x43, 0x09, 0x20, 0x38, 0x2D, 0x1A, 0x37,
	0x56, 0x33, 0x6D, 0x35, 0x2C, 0x57, 0x3D, 0x37, 0x2D, 0x52, 0x1A, 0x2C,
	0x72, 0x5D, 0x31, 0x3A, 0x1E, 0x69, 0x16, 0x3B, 0x04, 0x18, 0x7B, 0x2E,
	0x58, 0x1B, 0x11, 0x00, 0x59, 0x57, 0x5D, 0x18, 0x37, 0x3E, 0x08, 0x08,
	0x1F, 0x75, 0x2A, 0x0F, 0x00, 0x2E, 0x15, 0x0D, 0x31, 0x1F, 0x3F, 0x2C,
	0x05, 0x06, 0x01, 0x52, 0x37, 0x14, 0x59, 0x16, 0x1A, 0x0F, 0x54, 0x51,
	0x3A, 0x39, 0x7A, 0x16, 0x36, 0x25, 0x1D, 0x06, 0x29, 0x28, 0x20, 0x5A,
	0x0D, 0x01, 0x19, 0x04, 0x26, 0x04, 0x0E, 0x34, 0x0A, 0x0C, 0x18, 0x5D,
	0x31, 0x0A, 0x20, 0x72, 0x07, 0x59, 0x29, 0x1C, 0x06, 0x06, 0x58, 0x06,
	0x00, 0x03, 0x1E, 0x38, 0x0B, 0x04, 0x25, 0x3A, 0x24, 0x20, 0x25, 0x30,
	0x01, 0x24, 0x3F, 0x20, 0x72, 0x43, 0x2B, 0x24, 0x05, 0x13, 0x2E, 0x2E,
	0x21, 0x18, 0x1A, 0x00, 0x37, 0x22, 0x40, 0x11, 0x0E, 0x2F, 0x1C, 0x13,
	0x2B, 0x38, 0x27, 0x39, 0x53, 0x12, 0x03, 0x56, 0x5E, 0x25, 0x10, 0x18,
	0x55, 0x1D, 0x5B, 0x17, 0x1B, 0x12, 0x1C, 0x44, 0x01, 0x1E, 0x39, 0x22,
	0x19, 0x29, 0x07, 0x27, 0x22, 0x26, 0x35, 0x3F, 0x2D, 0x41, 0x53, 0x26,
	0x09, 0x2E, 0x45, 0x5E, 0x04, 0x5C, 0x2B, 0x5F, 0x44, 0x30, 0x3C, 0x52,
	0x20, 0x13, 0x07, 0x1E, 0x59, 0x0B, 0x44, 0x37, 0x3D, 0x27, 0x5A, 0x5B,
	0x0E, 0x3D, 0x2C, 0x3D, 0x3D, 0x30, 0x0F, 0x37, 0x1C, 0x2D, 0x05, 0x58,
	0x23, 0x1F, 0x11, 0x30, 0x0E, 0x59, 0x0D, 0x5F, 0x37, 0x5D, 0x30, 0x05,
	0x1F, 0x00, 0x27, 0x16, 0x0D, 0x29, 0x75, 0x20, 0x57, 0x29, 0x3C, 0x24,
	0x58, 0x24, 0x25, 0x33, 0x33, 0x09, 0x0D, 0x1E, 0x39, 0x06, 0x0E, 0x0E,
	0x07, 0x2F, 0x0E, 0x21, 0x26, 0x1B, 0x08, 0x77, 0x14, 0x37, 0x5D, 0x59,
	0x36, 0x26, 0x31, 0x3D, 0x20, 0x35, 0x5E, 0x17, 0x5A, 0x05, 0x29, 0x5F,
	0x57, 0x26, 0x33, 0x17, 0x20, 0x35, 0x41, 0x38, 0x70, 0x2E, 0x30, 0x07,
	0x3A, 0x09, 0x0A, 0x2B, 0x56, 0x2F, 0x32, 0x20, 0x2C, 0x56, 0x27, 0x2B,
	0x03, 0x30, 0x0F, 0x5D, 0x3A, 0x2A, 0x2A, 0x3D, 0x0A, 0x70, 0x1D, 0x33,
	0x5D, 0x25, 0x2D, 0x18, 0x36, 0x34, 0x1F, 0x0C, 0x2B, 0x25, 0x21, 0x04,
	0x08, 0x1F, 0x15, 0x2C, 0x38, 0x03, 0x0D, 0x32, 0x3E, 0x3A, 0x07, 0x0D,
	0x34, 0x37, 0x24, 0x16, 0x55, 0x2F, 0x09, 0x1E, 0x16, 0x22, 0x08, 0x2D,
	0x5E, 0x3B, 0x3C, 0x0A, 0x3B, 0x40, 0x2D, 0x06, 0x04, 0x1E, 0x19, 0x1B,
	0x1E, 0x03, 0x29, 0x2A, 0x2F, 0x47, 0x55, 0x3B, 0x2E, 0x36, 0x3C, 0x53,
	0x04, 0x32, 0x3B, 0x02, 0x31, 0x36, 0x13, 0x13, 0x3C, 0x26, 0x5C, 0x26,
	0x0A, 0x29, 0x12, 0x0C, 0x29, 0x16, 0x39, 0x36, 0x1D, 0x26, 0x05, 0x01,
	0x15, 0x5B, 0x33, 0x34, 0x38, 0x08, 0x34, 0x21, 0x75, 0x27, 0x0D, 0x23,
	0x1F, 0x76, 0x5E, 0x50, 0x37, 0x08, 0x15, 0x08, 0x03, 0x3E, 0x21, 0x09,
	0x06, 0x3B, 0x06, 0x26, 0x2C, 0x54, 0x53, 0x34, 0x53, 0x30, 0x38, 0x20,
	0x0A, 0x23, 0x7B, 0x27, 0x28, 0x0D, 0x32, 0x32, 0x28, 0x58, 0x5A, 0x1B,
	0x0F, 0x20, 0x53, 0x3D, 0x5A, 0x26, 0x04, 0x16, 0x1A, 0x20, 0x6D, 0x19,
	0x14, 0x28, 0x24, 0x2C, 0x06, 0x25, 0x2A, 0x5E, 0x29, 0x0B, 0x3B, 0x5F,
	0x1F, 0x06, 0x04, 0x0F, 0x2F, 0x5D, 0x23, 0x36, 0x2F, 0x0A, 0x40, 0x0F,
	0x25, 0x31, 0x21, 0x25, 0x0D, 0x5A, 0x0F, 0x03, 0x2D, 0x29, 0x47, 0x05,
	0x01, 0x3F, 0x7B, 0x21, 0x2A, 0x1F, 0x27, 0x1A, 0x1F, 0x18, 0x5E, 0x22,
	0x08, 0x02, 0x13, 0x5E, 0x5B, 0x0A, 0x2B, 0x4E, 0x37, 0x00, 0x2E, 0x00,
	0x17, 0x00, 0x0C, 0x2C, 0x3F, 0x09, 0x01, 0x08, 0x23, 0x38, 0x27, 0x5A,
	0x2D, 0x0E, 0x5A, 0x29, 0x02, 0x1F, 0x06, 0x01, 0x2C, 0x03, 0x06, 0x06,
	0x15, 0x09, 0x38, 0x06, 0x73, 0x59, 0x56, 0x23, 0x5E, 0x00, 0x01, 0x2F,
	0x3E, 0x5C, 0x1A, 0x26, 0x4A, 0x01, 0x03, 0x17, 0x00, 0x59, 0x14, 0x2C,
	0x33, 0x07, 0x20, 0x17, 0x5B, 0x75, 0x08, 0x25, 0x17, 0x0D, 0x33, 0x0B,
	0x55, 0x5E, 0x05, 0x15, 0x04, 0x57, 0x26, 0x02, 0x18, 0x24, 0x50, 0x09,
	0x20, 0x29, 0x5F, 0x36, 0x06, 0x5D, 0x33, 0x27, 0x3B, 0x26, 0x58, 0x35,
	0x1D, 0x0E, 0x2B, 0x23, 0x14, 0x39, 0x20, 0x2A, 0x2C, 0x0A, 0x2A, 0x59,
	0x34, 0x01, 0x75, 0x23, 0x28, 0x41, 0x3C, 0x11, 0x0E, 0x57, 0x2D, 0x1D,
	0x17, 0x38, 0x24, 0x57, 0x0F, 0x12, 0x24, 0x50, 0x1E, 0x26, 0x07, 0x1F,
	0x13, 0x45, 0x18, 0x2D, 0x2A, 0x33, 0x06, 0x5B, 0x2B, 0x27, 0x09, 0x37,
	0x44, 0x70, 0x05, 0x38, 0x07, 0x26, 0x26, 0x02, 0x11, 0x1C, 0x29, 0x2B,
	0x01, 0x08, 0x02, 0x02, 0x00, 0x3E, 0x29, 0x21, 0x1F, 0x75, 0x2D, 0x2B,
	0x2B, 0x1C, 0x05, 0x3C, 0x0B, 0x34, 0x20, 0x2D, 0x5D, 0x00, 0x20, 0x2D,
	0x7B, 0x2B, 0x09, 0x08, 0x11, 0x23, 0x3A, 0x0E, 0x0A, 0x04, 0x32, 0x3B,
	0x19, 0x58, 0x21, 0x77, 0x27, 0x27, 0x1F, 0x2A, 0x10, 0x3F, 0x15, 0x03,
	0x3E, 0x38, 0x1F, 0x58, 0x03, 0x18, 0x0A, 0x25, 0x0E, 0x1A, 0x3C, 0x38,
	0x0D, 0x22, 0x2D, 0x2D, 0x1A, 0x01, 0x36, 0x56, 0x33, 0x7A, 0x3C, 0x59,
	0x5E, 0x31, 0x2D, 0x47, 0x22, 0x58, 0x23, 0x09, 0x21, 0x36, 0x05, 0x58,
	0x6D, 0x20, 0x32, 0x37, 0x58, 0x2D, 0x23, 0x4E, 0x1A, 0x2D, 0x16, 0x0E,
	0x38, 0x1A, 0x04, 0x00, 0x06, 0x58, 0x05, 0x2C, 0x2E, 0x03, 0x09, 0x34,
	0x3F, 0x7A, 0x3F, 0x2D, 0x07, 0x0E, 0x03, 0x54, 0x09, 0x0D, 0x26, 0x70,
	0x28, 0x15, 0x1D, 0x5E, 0x75, 0x23, 0x27, 0x19, 0x26, 0x1B, 0x08, 0x2D,
	0x2F, 0x0A, 0x36, 0x43, 0x31, 0x0D, 0x0C, 0x29, 0x14, 0x23, 0x36, 0x3A,
	0x15, 0x3E, 0x15, 0x5E, 0x0A, 0x24, 0x3F, 0x22, 0x36, 0x07, 0x36, 0x3D,
	0x2E, 0x02, 0x31, 0x69, 0x27, 0x23, 0x03, 0x3C, 0x2B, 0x26, 0x13, 0x38,
	0x05, 0x09, 0x16, 0x31, 0x5B, 0x11, 0x03, 0x59, 0x19, 0x00, 0x2A, 0x34,
	0x39, 0x27, 0x0F, 0x21, 0x36, 0x16, 0x22, 0x21, 0x03, 0x1B, 0x28, 0x29,
	0x3F, 0x1D, 0x04, 0x1F, 0x23, 0x29, 0x09, 0x20, 0x05, 0x2C, 0x14, 0x24,
	0x3B, 0x23, 0x19, 0x2B, 0x5E, 0x2F, 0x2A, 0x0A, 0x26, 0x1F, 0x18, 0x07,
	0x33, 0x1D, 0x31, 0x00, 0x08, 0x34, 0x00, 0x13, 0x15, 0x03, 0x2B, 0x37,
	0x22, 0x07, 0x1E, 0x0C, 0x3F, 0x52, 0x71, 0x3A, 0x37, 0x1C, 0x29, 0x09,
	0x3B, 0x4E, 0x2B, 0x13, 0x14, 0x36, 0x0E, 0x36, 0x0D, 0x77, 0x3E, 0x2B,
	0x2D, 0x5D, 0x7B, 0x29, 0x20, 0x08, 0x38, 0x20, 0x06, 0x4A, 0x20, 0x5A,
	0x36, 0x43, 0x09, 0x04, 0x3D, 0x2C, 0x08, 0x2C, 0x01, 0x3E, 0x2C, 0x3F,
	0x04, 0x3D, 0x1E, 0x17, 0x1C, 0x31, 0x20, 0x3C, 0x0D, 0x29, 0x0F, 0x00,
	0x19, 0x17, 0x05, 0x32, 0x14, 0x07, 0x37, 0x2B, 0x26, 0x27, 0x0F, 0x23,
	0x08, 0x20, 0x58, 0x5A, 0x0B, 0x0E, 0x2E, 0x1A, 0x40, 0x35, 0x0E, 0x26,
	0x41, 0x02, 0x36, 0x36, 0x35, 0x39, 0x12, 0x2F, 0x28, 0x27, 0x26, 0x0E,
	0x06, 0x0E, 0x24, 0x1F, 0x02, 0x14, 0x0F, 0x20, 0x16, 0x18, 0x08, 0x23,
	0x0F, 0x3A, 0x3C, 0x18, 0x27, 0x31, 0x29, 0x27, 0x06, 0x3B, 0x19, 0x5C,
	0x24, 0x0C, 0x19, 0x25, 0x0D, 0x04, 0x25, 0x5A, 0x05, 0x0A, 0x32, 0x3B,
	0x21, 0x56, 0x5E, 0x25, 0x17, 0x0F, 0x29, 0x03, 0x3A, 0x76, 0x01, 0x36,
	0x39, 0x38, 0x25, 0x0B, 0x35, 0x2F, 0x23, 0x04, 0x39, 0x2D, 0x16, 0x07,
	0x0C, 0x0B, 0x10, 0x27, 0x3E, 0x0F, 0x2D, 0x18, 0x21, 0x1C, 0x07, 0x0E,
	0x02, 0x3C, 0x33, 0x77, 0x26, 0x50, 0x29, 0x3F, 0x34, 0x5E, 0x27, 0x07,
	0x29, 0x7B, 0x3C, 0x25, 0x1E, 0x01, 0x32, 0x1B, 0x04, 0x5E, 0x11, 0x31,
	0x2E, 0x2B, 0x03, 0x5F, 0x0B, 0x09, 0x0D, 0x3A, 0x39, 0x71, 0x18, 0x31,
	0x3E, 0x31, 0x0E, 0x5D, 0x0E, 0x56, 0x04, 0x25, 0x20, 0x37, 0x2A, 0x21,
	0x0C, 0x3B, 0x1B, 0x0F, 0x06, 0x0A, 0x3C, 0x06, 0x57, 0x1C, 0x09, 0x5B,
	0x10, 0x34, 0x0D, 0x29, 0x06, 0x58, 0x5E, 0x2E, 0x70, 0x09, 0x1B, 0x39,
	0x1B, 0x21, 0x09, 0x13, 0x1A, 0x11, 0x0D, 0x2A, 0x20, 0x18, 0x08, 0x34,
	0x27, 0x37, 0x39, 0x04, 0x30, 0x15, 0x15, 0x37, 0x38, 0x71, 0x04, 0x2C,
	0x04, 0x24, 0x13, 0x3C, 0x0B, 0x23, 0x3A, 0x31, 0x5D, 0x39, 0x08, 0x53,
	0x0E, 0x0E, 0x28, 0x1E, 0x24, 0x2C, 0x3F, 0x0E, 0x2D, 0x0F, 0x7A, 0x3B,
	0x57, 0x5C, 0x52, 0x1A, 0x5F, 0x38, 0x5B, 0x12, 0x0B, 0x39, 0x52, 0x18,
	0x44, 0x74, 0x3A, 0x57, 0x0F, 0x24, 0x1A, 0x18, 0x35, 0x2D, 0x5E, 0x21,
	0x1D, 0x38, 0x0A, 0x33, 0x74, 0x23, 0x24, 0x3E, 0x58, 0x7A, 0x5B, 0x24,
	0x39, 0x0C, 0x70, 0x24, 0x00, 0x14, 0x07, 0x21, 0x14, 0x4A, 0x2B, 0x2A,
	0x2A, 0x5C, 0x2C, 0x24, 0x2C, 0x01, 0x0A, 0x24, 0x1A, 0x03, 0x10, 0x08,
	0x07, 0x21, 0x19, 0x2A, 0x28, 0x4A, 0x06, 0x5B, 0x07, 0x3D, 0x55, 0x0C,
	0x3E, 0x25, 0x36, 0x08, 0x23, 0x5F, 0x21, 0x18, 0x2A, 0x0A, 0x01, 0x69,
	0x2E, 0x4E, 0x3A, 0x2D, 0x08, 0x1B, 0x20, 0x20, 0x13, 0x26, 0x07, 0x57,
	0x41, 0x52, 0x36, 0x22, 0x2C, 0x39, 0x2D, 0x28, 0x5C, 0x17, 0x02, 0x2A,
	0x30, 0x58, 0x2D, 0x5F, 0x3D, 0x05, 0x03, 0x19, 0x07, 0x11, 0x15, 0x16,
	0x39, 0x1A, 0x21, 0x73, 0x3A, 0x2C, 0x3D, 0x5F, 0x2C, 0x27, 0x0A, 0x5F,
	0x21, 0x21, 0x05, 0x3B, 0x21, 0x0C, 0x0E, 0x2A, 0x2F, 0x01, 0x04, 0x20,
	0x21, 0x22, 0x3B, 0x5B, 0x27, 0x1F, 0x08, 0x3B, 0x5B, 0x01, 0x3C, 0x22,
	0x22, 0x22, 0x04, 0x05, 0x2B, 0x1D, 0x03, 0x18, 0x2D, 0x10, 0x39, 0x3E,
	0x03, 0x26, 0x3B, 0x2D, 0x5C, 0x3A, 0x3F, 0x34, 0x06, 0x1B, 0x2E, 0x1B,
	0x07, 0x3B, 0x59, 0x0F, 0x36, 0x32, 0x5C, 0x2E, 0x23, 0x55, 0x0B, 0x19,
	0x40, 0x2B, 0x1B, 0x03, 0x36, 0x07, 0x7B, 0x00, 0x16, 0x5C, 0x18, 0x36,
	0x2B, 0x50, 0x59, 0x19, 0x35, 0x55, 0x32, 0x06, 0x0A, 0x36, 0x06, 0x16,
	0x03, 0x1D, 0x12, 0x3F, 0x0A, 0x17, 0x3A, 0x76, 0x38, 0x38, 0x41, 0x26,
	0x2B, 0x34, 0x31, 0x2A, 0x5F, 0x77, 0x3A, 0x57, 0x3A, 0x3D, 0x6D, 0x2E,
	0x00, 0x03, 0x01, 0x3A, 0x02, 0x2C, 0x3C, 0x59, 0x06, 0x19, 0x14, 0x06,
	0x28, 0x73, 0x0B, 0x24, 0x23, 0x52, 0x15, 0x5D, 0x29, 0x00, 0x09, 0x12,
	0x24, 0x2F, 0x0C, 0x59, 0x04, 0x47, 0x14, 0x5E, 0x03, 0x2B, 0x18, 0x3B,
	0x45, 0x25, 0x35, 0x59, 0x04, 0x1E, 0x5A, 0x38, 0x5E, 0x2C, 0x24, 0x03,
	0x05, 0x58, 0x07, 0x1A, 0x23, 0x12, 0x36, 0x16, 0x1B, 0x21, 0x28, 0x28,
	0x11, 0x3C, 0x12, 0x37, 0x58, 0x29, 0x2F, 0x25, 0x2A, 0x5E, 0x12, 0x5B,
	0x33, 0x0F, 0x0A, 0x09, 0x2F, 0x22, 0x26, 0x28, 0x29, 0x2F, 0x5E, 0x38,
	0x23, 0x2C, 0x24, 0x03, 0x25, 0x58, 0x51, 0x1C, 0x3B, 0x76, 0x0F, 0x15,
	0x26, 0x27, 0x18, 0x14, 0x53, 0x23, 0x5E, 0x2A, 0x28, 0x55, 0x0B, 0x27,
	0x0D, 0x3A, 0x1B, 0x25, 0x5F, 0x13, 0x03, 0x2E, 0x5F, 0x58, 0x01, 0x58,
	0x0D, 0x1D, 0x25, 0x73, 0x24, 0x20, 0x5B, 0x1C, 0x0D, 0x21, 0x35, 0x06,
	0x26, 0x0B, 0x0F, 0x0B, 0x26, 0x2F, 0x20, 0x07, 0x02, 0x0B, 0x33, 0x2C,
	0x1F, 0x28, 0x36, 0x2F, 0x0C, 0x0B, 0x56, 0x0C, 0x24, 0x27, 0x16, 0x09,
	0x0D, 0x2F, 0x05, 0x24, 0x32, 0x14, 0x07, 0x21, 0x1B, 0x04, 0x2B, 0x0A,
	0x06, 0x18, 0x05, 0x17, 0x1E, 0x0B, 0x5B, 0x25, 0x2F, 0x3A, 0x74, 0x24,
	0x2E, 0x2C, 0x11, 0x2F, 0x0F, 0x28, 0x3A, 0x2F, 0x2A, 0x1D, 0x14, 0x5A,
	0x53, 0x2C, 0x3C, 0x38, 0x19, 0x06, 0x07, 0x0E, 0x09, 0x45, 0x5B, 0x21,
	0x55, 0x0F, 0x2D, 0x5F, 0x2F, 0x21, 0x2E, 0x02, 0x23, 0x09, 0x5B, 0x06,
	0x0D, 0x2A, 0x70, 0x24, 0x00, 0x14, 0x07, 0x21, 0x14, 0x4A, 0x2B, 0x2A,
	0x2A, 0x5C, 0x2C, 0x0D, 0x2F, 0x2C, 0x21, 0x55, 0x19, 0x06, 0x0A, 0x28,
	0x1B, 0x59, 0x01, 0x3B, 0x0F, 0x58, 0x04, 0x28, 0x1B, 0x3E, 0x14, 0x26,
	0x5C, 0x10, 0x16, 0x53, 0x0D, 0x27, 0x2B, 0x35, 0x16, 0x58, 0x3E, 0x21,
	0x1E, 0x14, 0x2C, 0x1C, 0x06, 0x35, 0x05, 0x1C, 0x24, 0x14, 0x16, 0x29,
	0x5A, 0x3A, 0x01, 0x24, 0x30, 0x16, 0x1C, 0x0D, 0x0F, 0x1B, 0x04, 0x28,
	0x1B, 0x0F, 0x31, 0x38, 0x33, 0x12, 0x07, 0x54, 0x0C, 0x24, 0x05, 0x1B,
	0x0B, 0x0D, 0x25, 0x70, 0x28, 0x0F, 0x1D, 0x5F, 0x1A, 0x21, 0x1B, 0x06,
	0x3E, 0x25, 0x59, 0x39, 0x0D, 0x27, 0x2B, 0x2B, 0x16, 0x59, 0x3E, 0x21,
	0x1E, 0x14, 0x20, 0x1C, 0x25, 0x21, 0x2C, 0x06, 0x2F, 0x2D, 0x0F, 0x54,
	0x26, 0x24, 0x05, 0x1B, 0x38, 0x3C, 0x21, 0x1A, 0x0A, 0x06, 0x5B, 0x09,
	0x0D, 0x2B, 0x1B, 0x04, 0x18, 0x08, 0x5F, 0x25, 0x26, 0x0C, 0x76, 0x34,
	0x02, 0x59, 0x02, 0x17, 0x1B, 0x19, 0x3B, 0x08, 0x30, 0x19, 0x27, 0x19,
	0x27, 0x1B, 0x0A, 0x13, 0x21, 0x29, 0x38, 0x0B, 0x02, 0x27, 0x01, 0x06,
	0x35, 0x30, 0x5B, 0x23, 0x0D, 0x2B, 0x1B, 0x5A, 0x23, 0x74, 0x5B, 0x59,
	0x26, 0x27, 0x18, 0x1B, 0x53, 0x23, 0x31, 0x2A, 0x23, 0x55, 0x0D, 0x52,
	0x0A, 0x2F, 0x56, 0x03, 0x08, 0x01, 0x01, 0x29, 0x25, 0x11, 0x2A, 0x0F,
	0x16, 0x45, 0x2D, 0x23, 0x28, 0x15, 0x0A, 0x13, 0x0D, 0x21, 0x25, 0x06,
	0x2E, 0x0B, 0x0A, 0x25, 0x26, 0x22, 0x77, 0x1B, 0x53, 0x3E, 0x29, 0x38,
	0x1E, 0x17, 0x19, 0x08, 0x36, 0x02, 0x25, 0x37, 0x13, 0x2F, 0x29, 0x56,
	0x06, 0x11, 0x72, 0x0F, 0x2D, 0x1B, 0x31, 0x35, 0x27, 0x38, 0x0D, 0x19,
	0x0D, 0x2A, 0x1B, 0x2A, 0x5F, 0x14, 0x03, 0x2E, 0x5F, 0x58, 0x07, 0x58,
	0x16, 0x21, 0x2E, 0x13, 0x04, 0x59, 0x23, 0x08, 0x28, 0x02, 0x25, 0x37,
	0x26, 0x08, 0x07, 0x13, 0x3E, 0x5F, 0x21, 0x18, 0x29, 0x22, 0x31, 0x3A,
	0x5E, 0x2C, 0x5B, 0x03, 0x06, 0x58, 0x04, 0x22, 0x24, 0x14, 0x16, 0x2A,
	0x5A, 0x3A, 0x2D, 0x23, 0x50, 0x5D, 0x28, 0x76, 0x00, 0x12, 0x20, 0x5A,
	0x0A, 0x2D, 0x54, 0x19, 0x24, 0x0F, 0x38, 0x09, 0x23, 0x22, 0x21, 0x06,
	0x29, 0x2A, 0x09, 0x29, 0x0F, 0x4A, 0x36, 0x05, 0x31, 0x25, 0x39, 0x2A,
	0x25, 0x25, 0x5B, 0x03, 0x21, 0x0E, 0x38, 0x04, 0x02, 0x2A, 0x2C, 0x0A,
	0x3F, 0x1B, 0x02, 0x08, 0x35, 0x09, 0x24, 0x0F, 0x2F, 0x36, 0x08, 0x18,
	0x1B, 0x22, 0x75, 0x28, 0x20, 0x3F, 0x5D, 0x0A, 0x23, 0x23, 0x14, 0x06,
	0x21, 0x25, 0x35, 0x2A, 0x03, 0x2F, 0x19, 0x55, 0x56, 0x05, 0x12, 0x35,
	0x16, 0x03, 0x2E, 0x20, 0x04, 0x4A, 0x5E, 0x08, 0x7B, 0x02, 0x22, 0x5A,
	0x06, 0x0F, 0x23, 0x0D, 0x26, 0x20, 0x75, 0x0B, 0x02, 0x2F, 0x59, 0x0A,
	0x0D, 0x1B, 0x02, 0x08, 0x3A, 0x47, 0x24, 0x2F, 0x03, 0x72, 0x21, 0x02,
	0x2A, 0x05, 0x0F, 0x58, 0x16, 0x03, 0x23, 0x06, 0x18, 0x37, 0x14, 0x5E,
	0x0D, 0x3B, 0x1B, 0x06, 0x18, 0x0B, 0x5F, 0x25, 0x0A, 0x0C, 0x77, 0x5B,
	0x2E, 0x28, 0x11, 0x0F, 0x58, 0x37, 0x27, 0x24, 0x14, 0x5F, 0x22, 0x5A,
	0x03, 0x31, 0x23, 0x50, 0x26, 0x20, 0x75, 0x06, 0x02, 0x27, 0x2F, 0x06,
	0x25, 0x30, 0x58, 0x23, 0x0D, 0x3E, 0x1B, 0x06, 0x18, 0x05, 0x29, 0x2A,
	0x38, 0x58, 0x76, 0x23, 0x36, 0x14, 0x03, 0x31, 0x58, 0x56, 0x2D, 0x0F,
	0x35, 0x14, 0x55, 0x21, 0x2D, 0x71, 0x23, 0x55, 0x02, 0x26, 0x0F, 0x3A,
	0x29, 0x25, 0x5C, 0x2A, 0x0F, 0x22, 0x5C, 0x23, 0x74, 0x16, 0x06, 0x0D,
	0x5F, 0x0A, 0x2F, 0x28, 0x19, 0x59, 0x07, 0x23, 0x33, 0x14, 0x02, 0x0F,
	0x24, 0x0F, 0x37, 0x2C, 0x2E, 0x26, 0x4E, 0x2A, 0x2D, 0x25, 0x5B, 0x03,
	0x21, 0x2C, 0x38, 0x02, 0x12, 0x27, 0x0D, 0x06, 0x14, 0x33, 0x19, 0x1E,
	0x77, 0x34, 0x20, 0x28, 0x03, 0x70, 0x1F, 0x55, 0x36, 0x26, 0x34, 0x04,
	0x2E, 0x09, 0x5F, 0x0A, 0x23, 0x23, 0x14, 0x02, 0x21, 0x26, 0x0B, 0x2A,
	0x2E, 0x13, 0x58, 0x03, 0x1C, 0x1E, 0x12, 0x27, 0x1B, 0x5C, 0x2E, 0x0E,
	0x04, 0x53, 0x5E, 0x08, 0x36, 0x02, 0x31, 0x37, 0x1C, 0x69, 0x2A, 0x08,
	0x2A, 0x1B, 0x26, 0x15, 0x14, 0x27, 0x27, 0x06, 0x22, 0x33, 0x17, 0x1E,
	0x77, 0x34, 0x20, 0x0A, 0x03, 0x35, 0x21, 0x02, 0x2A, 0x05, 0x07, 0x58,
	0x1B, 0x21, 0x2E, 0x0B, 0x04, 0x16, 0x5D, 0x33, 0x21, 0x47, 0x39, 0x00,
	0x18, 0x0B, 0x34, 0x25, 0x20, 0x0C, 0x75, 0x0E, 0x2E, 0x0B, 0x11, 0x2A,
	0x0F, 0x25, 0x29, 0x23, 0x11, 0x16, 0x0D, 0x0D, 0x1C, 0x27, 0x29, 0x00,
	0x2A, 0x1F, 0x26, 0x15, 0x14, 0x27, 0x5C, 0x06, 0x2D, 0x30, 0x58, 0x23,
	0x0D, 0x2E, 0x1B, 0x03, 0x08, 0x0B, 0x38, 0x25, 0x2C, 0x01, 0x36, 0x34,
	0x07, 0x09, 0x5E, 0x20, 0x23, 0x26, 0x14, 0x01, 0x31, 0x26, 0x52, 0x2A,
	0x23, 0x25, 0x58, 0x39, 0x0D, 0x5C, 0x2B, 0x39, 0x16, 0x16, 0x3E, 0x21,
	0x1E, 0x14, 0x28, 0x1C, 0x0E, 0x35, 0x07, 0x1C, 0x24, 0x00, 0x16, 0x06,
	0x0D, 0x22, 0x28, 0x28, 0x38, 0x3F, 0x5E, 0x0A, 0x23, 0x26, 0x16, 0x1C,
	0x21, 0x23, 0x39, 0x00, 0x18, 0x0B, 0x34, 0x25, 0x20, 0x0C, 0x75, 0x0E,
	0x2E, 0x0B, 0x11, 0x2A, 0x0F, 0x25, 0x29, 0x23, 0x11, 0x16, 0x0D, 0x0D,
	0x1C, 0x27, 0x29, 0x00, 0x2A, 0x1F, 0x26, 0x15, 0x14, 0x27, 0x5C, 0x06,
	0x2D, 0x30, 0x58, 0x23, 0x0D, 0x2E, 0x1B, 0x03, 0x08, 0x0B, 0x38, 0x25,
	0x06, 0x06, 0x2E, 0x0F, 0x4A, 0x3A, 0x07, 0x31, 0x58, 0x03, 0x2D, 0x25,
	0x35, 0x5F, 0x38, 0x21, 0x0E, 0x38, 0x04, 0x02, 0x14, 0x24, 0x04, 0x3F,
	0x25, 0x02, 0x0F, 0x35, 0x19, 0x28, 0x0C, 0x2F, 0x36, 0x3E, 0x18, 0x1B,
	0x5F, 0x71, 0x2F, 0x20, 0x19, 0x12, 0x07, 0x23, 0x09, 0x14, 0x00, 0x21,
	0x58, 0x03, 0x2C, 0x03, 0x0D, 0x00, 0x05, 0x45, 0x2F, 0x2E, 0x1A, 0x30,
	0x19, 0x26, 0x06, 0x15, 0x24, 0x38, 0x1F, 0x38, 0x06, 0x32, 0x5E, 0x58,
	0x04, 0x1F, 0x59, 0x5B, 0x5A, 0x3A, 0x20, 0x52, 0x45, 0x24, 0x2C, 0x55,
	0x32, 0x57, 0x12, 0x76, 0x21, 0x22, 0x18, 0x21, 0x0C, 0x0E, 0x2E, 0x14,
	0x0A, 0x13, 0x34, 0x35, 0x41, 0x27, 0x34, 0x29, 0x2B, 0x0B, 0x5D, 0x23,
	0x07, 0x30, 0x34, 0x2F, 0x25, 0x5D, 0x52, 0x08, 0x1B, 0x00, 0x1F, 0x52,
	0x24, 0x5C, 0x74, 0x03, 0x53, 0x36, 0x18, 0x20, 0x3B, 0x4A, 0x22, 0x2C,
	0x7B, 0x5D, 0x35, 0x5E, 0x00, 0x1B, 0x14, 0x0A, 0x58, 0x29, 0x3A, 0x0F,
	0x52, 0x2A, 0x3F, 0x30, 0x2F, 0x54, 0x34, 0x5A, 0x27, 0x01, 0x0B, 0x29,
	0x05, 0x12, 0x5B, 0x27, 0x14, 0x32, 0x03, 0x09, 0x0D, 0x04, 0x0A, 0x0A,
	0x20, 0x36, 0x59, 0x24, 0x72, 0x2B, 0x52, 0x3C, 0x3A, 0x2C, 0x1D, 0x55,
	0x27, 0x3D, 0x1B, 0x36, 0x29, 0x27, 0x5E, 0x35, 0x5E, 0x25, 0x2C, 0x1A,
	0x0B, 0x28, 0x3B, 0x14, 0x59, 0x0F, 0x26, 0x09, 0x29, 0x5F, 0x24, 0x18,
	0x29, 0x3E, 0x31, 0x35, 0x19, 0x2B, 0x04, 0x2F, 0x32, 0x3E, 0x18, 0x1B,
	0x5F, 0x0A, 0x2D, 0x2F, 0x06, 0x59, 0x31, 0x59, 0x39, 0x23, 0x0D, 0x2A,
	0x2D, 0x28, 0x0A, 0x2F, 0x0A, 0x2D, 0x54, 0x14, 0x24, 0x0F, 0x26, 0x09,
	0x19, 0x5B, 0x14, 0x0F, 0x4A, 0x3A, 0x07, 0x31, 0x58, 0x03, 0x2D, 0x25,
	0x35, 0x5F, 0x38, 0x21, 0x0E, 0x38, 0x04, 0x02, 0x14, 0x24, 0x04, 0x3F,
	0x25, 0x02, 0x0F, 0x35, 0x19, 0x28, 0x0C, 0x2F, 0x36, 0x3E, 0x18, 0x1B,
	0x5F, 0x71, 0x2F, 0x20, 0x19, 0x12, 0x07, 0x23, 0x09, 0x14, 0x00, 0x21,
	0x58, 0x03, 0x2A, 0x03, 0x1B, 0x1D, 0x56, 0x56, 0x23, 0x0E, 0x36, 0x16,
	0x5C, 0x26, 0x18, 0x04, 0x2E, 0x5A, 0x08, 0x7B, 0x24, 0x22, 0x59, 0x06,
	0x21, 0x2F, 0x0C, 0x26, 0x20, 0x38, 0x04, 0x02, 0x19, 0x40, 0x04, 0x0D,
	0x25, 0x1A, 0x0F, 0x3A, 0x23, 0x2C, 0x2A, 0x03, 0x07, 0x25, 0x07, 0x2A,
	0x23, 0x0B, 0x59, 0x16, 0x29, 0x24, 0x71, 0x3E, 0x23, 0x1E, 0x38, 0x24,
	0x1B, 0x19, 0x37, 0x24, 0x70, 0x16, 0x09, 0x1D, 0x5E, 0x75, 0x2F, 0x29,
	0x19, 0x53, 0x17, 0x0F, 0x2D, 0x1B, 0x3D, 0x35, 0x2E, 0x38, 0x0A, 0x19,
	0x0D, 0x2A, 0x1B, 0x22, 0x5F, 0x16, 0x03, 0x2E, 0x2C, 0x11, 0x25, 0x0F,
	0x55, 0x00, 0x28, 0x1B, 0x1B, 0x19, 0x2B, 0x24, 0x05, 0x5C, 0x3B, 0x14,
	0x5E, 0x27, 0x09, 0x16, 0x06, 0x08, 0x0F, 0x5E, 0x25, 0x1A, 0x18, 0x77,
	0x5B, 0x2E, 0x28, 0x1C, 0x0F, 0x35, 0x05, 0x22, 0x24, 0x14, 0x16, 0x23,
	0x5A, 0x39, 0x2D, 0x23, 0x50, 0x5D, 0x20, 0x76, 0x06, 0x12, 0x23, 0x29,
	0x06, 0x03, 0x02, 0x5A, 0x23, 0x0D, 0x36, 0x16, 0x06, 0x26, 0x0D, 0x2B,
	0x2C, 0x38, 0x11, 0x77, 0x23, 0x36, 0x14, 0x03, 0x31, 0x25, 0x52, 0x2A,
	0x0F, 0x25, 0x59, 0x56, 0x21, 0x2D, 0x38, 0x21, 0x55, 0x38, 0x22, 0x0D,
	0x3A, 0x52, 0x2D, 0x5F, 0x2A, 0x1F, 0x2E, 0x5F, 0x23, 0x09, 0x5B, 0x0B,
	0x0D, 0x22, 0x06, 0x28, 0x28, 0x3F, 0x5D, 0x0A, 0x23, 0x33, 0x14, 0x03,
	0x31, 0x2B, 0x24, 0x1D, 0x3D, 0x71, 0x58, 0x2E, 0x39, 0x11, 0x2A, 0x1F,
	0x55, 0x59, 0x28, 0x26, 0x1B, 0x19, 0x5A, 0x24, 0x04, 0x5F, 0x2E, 0x5A,
	0x07, 0x0F, 0x21, 0x37, 0x26, 0x20, 0x75, 0x04, 0x02, 0x2D, 0x59, 0x0A,
	0x5A, 0x1B, 0x09, 0x08, 0x76, 0x24, 0x22, 0x27, 0x1C, 0x70, 0x29, 0x2E,
	0x3C, 0x11, 0x2A, 0x1F, 0x18, 0x21, 0x33, 0x09, 0x16, 0x53, 0x2B, 0x27,
	0x2A, 0x5E, 0x51, 0x0D, 0x1F, 0x2C, 0x3C, 0x38, 0x19, 0x40, 0x04, 0x05,
	0x25, 0x1E, 0x0F, 0x3B, 0x19, 0x28, 0x22, 0x2F, 0x0C, 0x3E, 0x18, 0x1B,
	0x5E, 0x1A, 0x2D, 0x05, 0x06, 0x1C, 0x0F, 0x0F, 0x25, 0x00, 0x2E, 0x76,
	0x16, 0x2E, 0x2B, 0x22, 0x2A, 0x1B, 0x52, 0x04, 0x1E, 0x12, 0x26, 0x1B,
	0x5C, 0x26, 0x08, 0x04, 0x26, 0x5A, 0x0D, 0x36, 0x24, 0x31, 0x34, 0x1C,
	0x37, 0x26, 0x0B, 0x2A, 0x1B, 0x10, 0x15, 0x14, 0x5A, 0x23, 0x03, 0x22,
	0x09, 0x5C, 0x18, 0x77, 0x34, 0x2C, 0x08, 0x03, 0x03, 0x25, 0x05, 0x2A,
	0x23, 0x03, 0x59, 0x1B, 0x21, 0x26, 0x08, 0x04, 0x16, 0x17, 0x3D, 0x21,
	0x47, 0x35, 0x02, 0x18, 0x76, 0x0E, 0x22, 0x20, 0x1C, 0x71, 0x35, 0x2E,
	0x0B, 0x11, 0x2A, 0x0F, 0x1B, 0x21, 0x2D, 0x11, 0x28, 0x0D, 0x0A, 0x1C,
	0x37, 0x25, 0x03, 0x2A, 0x1F, 0x10, 0x15, 0x14, 0x5A, 0x58, 0x01, 0x2D,
	0x16, 0x17, 0x2E, 0x0D, 0x04, 0x1B, 0x05, 0x08, 0x76, 0x0E, 0x25, 0x06,
	0x3E, 0x33, 0x5B, 0x59, 0x26, 0x27, 0x18, 0x1B, 0x53, 0x23, 0x31, 0x2A,
	0x23, 0x55, 0x0D, 0x52, 0x0A, 0x2F, 0x56, 0x03, 0x08, 0x01, 0x01, 0x29,
	0x25, 0x11, 0x2A, 0x0F, 0x16, 0x45, 0x2D, 0x23, 0x28, 0x15, 0x0A, 0x13,
	0x0D, 0x21, 0x25, 0x06, 0x2E, 0x0B, 0x0A, 0x25, 0x26, 0x22, 0x77, 0x1B,
	0x53, 0x2A, 0x28, 0x27, 0x27, 0x1B, 0x45, 0x23, 0x0E, 0x3E, 0x18, 0x5C,
	0x08, 0x26, 0x06, 0x2E, 0x37, 0x3A, 0x69, 0x24, 0x08, 0x14, 0x07, 0x21,
	0x15, 0x14, 0x2B, 0x20, 0x06, 0x18, 0x05, 0x19, 0x1E, 0x08, 0x0E, 0x25,
	0x0A, 0x39, 0x35, 0x23, 0x02, 0x2A, 0x01, 0x07, 0x58, 0x35, 0x2D, 0x23,
	0x0B, 0x14, 0x16, 0x5C, 0x3C, 0x0E, 0x02, 0x18, 0x0D, 0x52, 0x28, 0x2F,
	0x38, 0x3C, 0x1E, 0x0A, 0x5B, 0x33, 0x14, 0x59, 0x21, 0x20, 0x08, 0x37,
	0x1C, 0x74, 0x39, 0x02, 0x1C, 0x1E, 0x00, 0x1B, 0x25, 0x37, 0x0F, 0x30,
	0x23, 0x37, 0x14, 0x23, 0x76, 0x3D, 0x22, 0x26, 0x3A, 0x3A, 0x1B, 0x2E,
	0x0D, 0x11, 0x28, 0x2F, 0x38, 0x0D, 0x25, 0x2E, 0x34, 0x31, 0x05, 0x5E,
	0x20, 0x23, 0x26, 0x19, 0x01, 0x21, 0x22, 0x53, 0x2A, 0x05, 0x31, 0x58,
	0x39, 0x23, 0x11, 0x2A, 0x39, 0x06, 0x5B, 0x33, 0x21, 0x20, 0x08, 0x29,
	0x1C, 0x75, 0x39, 0x02, 0x1C, 0x1E, 0x0C, 0x1B, 0x06, 0x23, 0x26, 0x2A,
	0x28, 0x0E, 0x0D, 0x5E, 0x0A, 0x23, 0x26, 0x19, 0x5F, 0x1A, 0x27, 0x14,
	0x41, 0x29, 0x3B, 0x5E, 0x02, 0x20, 0x01, 0x05, 0x35, 0x35, 0x1B, 0x23,
	0x12, 0x3E, 0x16, 0x1B, 0x5E, 0x2C, 0x2D, 0x11, 0x06, 0x12, 0x31, 0x58,
	0x39, 0x23, 0x3B, 0x2A, 0x3B, 0x06, 0x59, 0x33, 0x21, 0x38, 0x0B, 0x2F,
	0x5F, 0x10, 0x2F, 0x29, 0x19, 0x13, 0x3B, 0x23, 0x02, 0x20, 0x0C, 0x35,
	0x0B, 0x32, 0x1D, 0x44, 0x2A, 0x15, 0x51, 0x0D, 0x1F, 0x2C, 0x24, 0x38,
	0x14, 0x06, 0x07, 0x3C, 0x09, 0x5A, 0x18, 0x77, 0x34, 0x2C, 0x1C, 0x03,
	0x01, 0x0B, 0x56, 0x36, 0x08, 0x0E, 0x05, 0x36, 0x19, 0x58, 0x17, 0x0F,
	0x25, 0x00, 0x2A, 0x76, 0x14, 0x2E, 0x2B, 0x1C, 0x2A, 0x15, 0x2C, 0x0D,
	0x25, 0x29, 0x16, 0x0A, 0x17, 0x18, 0x7B, 0x04, 0x22, 0x5A, 0x0F, 0x36,
	0x24, 0x2D, 0x34, 0x11, 0x70, 0x21, 0x31, 0x06, 0x32, 0x25, 0x5A, 0x39,
	0x0D, 0x19, 0x2B, 0x2F, 0x16, 0x14, 0x3E, 0x21, 0x1E, 0x14, 0x38, 0x1C,
	0x0A, 0x35, 0x02, 0x2A, 0x23, 0x03, 0x59, 0x19, 0x21, 0x26, 0x38, 0x04,
	0x22, 0x27, 0x08, 0x0C, 0x3A, 0x52, 0x2A, 0x07, 0x77, 0x5B, 0x22, 0x28,
	0x1C, 0x38, 0x35, 0x2E, 0x5C, 0x11, 0x2C, 0x1F, 0x55, 0x36, 0x2A, 0x3A,
	0x04, 0x51, 0x1D, 0x5E, 0x1A, 0x21, 0x29, 0x06, 0x2C, 0x25, 0x5B, 0x39,
	0x0D, 0x19, 0x2B, 0x23, 0x16, 0x19, 0x23, 0x03, 0x5A, 0x15, 0x24, 0x58,
	0x70, 0x2B, 0x28, 0x38, 0x27, 0x2B, 0x23, 0x05, 0x18, 0x3E, 0x28, 0x3A,
	0x04, 0x05, 0x33, 0x6D, 0x25, 0x09, 0x39, 0x1E, 0x13, 0x39, 0x0D, 0x17,
	0x11, 0x27, 0x3F, 0x09, 0x1A, 0x2E, 0x2A, 0x5D, 0x16, 0x41, 0x11, 0x1B,
	0x25, 0x11, 0x39, 0x40, 0x0A, 0x1E, 0x39, 0x1E, 0x25, 0x31, 0x2B, 0x06,
	0x45, 0x52, 0x27, 0x0A, 0x58, 0x21, 0x0D, 0x21, 0x5E, 0x23, 0x1F, 0x3E,
	0x32, 0x29, 0x19, 0x57, 0x3B, 0x2E, 0x09, 0x28, 0x00, 0x1C, 0x34, 0x26,
	0x2B, 0x3A, 0x1D, 0x72, 0x05, 0x04, 0x45, 0x52, 0x25, 0x1F, 0x02, 0x1D,
	0x0F, 0x72, 0x5F, 0x22, 0x36, 0x44, 0x1A, 0x01, 0x2F, 0x41, 0x3C, 0x75,
	0x21, 0x05, 0x09, 0x31, 0x07, 0x0A, 0x0C, 0x1A, 0x33, 0x07, 0x54, 0x2A,
	0x1E, 0x33, 0x08, 0x5B, 0x2D, 0x04, 0x1E, 0x2A, 0x34, 0x24, 0x28, 0x1C,
	0x74, 0x01, 0x18, 0x2F, 0x5D, 0x07, 0x5C, 0x56, 0x09, 0x28, 0x16, 0x2A,
	0x0B, 0x21, 0x39, 0x23, 0x28, 0x23, 0x23, 0x33, 0x17, 0x00, 0x20, 0x1E,
	0x28, 0x75, 0x1D, 0x22, 0x37, 0x19, 0x70, 0x3A, 0x36, 0x56, 0x3B, 0x25,
	0x23, 0x25, 0x5C, 0x39, 0x15, 0x1C, 0x03, 0x27, 0x29, 0x24, 0x1E, 0x03,
	0x21, 0x1D, 0x1B, 0x5E, 0x24, 0x17, 0x2C, 0x75, 0x5A, 0x27, 0x29, 0x38,
	0x16, 0x38, 0x31, 0x36, 0x04, 0x3B, 0x5E, 0x14, 0x58, 0x32, 0x37, 0x14,
	0x2D, 0x2B, 0x1A, 0x03, 0x3E, 0x35, 0x05, 0x53, 0x2E, 0x07, 0x34, 0x24,
	0x18, 0x11, 0x06, 0x09, 0x1D, 0x08, 0x3A, 0x21, 0x51, 0x5E, 0x5E, 0x71,
	0x3A, 0x54, 0x02, 0x59, 0x38, 0x2B, 0x03, 0x2B, 0x32, 0x17, 0x0D, 0x59,
	0x38, 0x38, 0x27, 0x23, 0x2C, 0x21, 0x22, 0x05, 0x3C, 0x32, 0x02, 0x2F,
	0x09, 0x1E, 0x50, 0x57, 0x33, 0x1A, 0x55, 0x13, 0x24, 0x01, 0x28, 0x1C,
	0x2D, 0x5C, 0x24, 0x3A, 0x25, 0x34, 0x14, 0x03, 0x2E, 0x58, 0x53, 0x3B,
	0x04, 0x32, 0x3F, 0x08, 0x00, 0x13, 0x38, 0x3A, 0x07, 0x45, 0x0D, 0x30,
	0x1A, 0x59, 0x18, 0x5B, 0x1A, 0x59, 0x4E, 0x45, 0x40, 0x74, 0x16, 0x4A,
	0x45, 0x5D, 0x30, 0x47, 0x36, 0x58, 0x44, 0x6D, 0x18, 0x14, 0x1F, 0x44,
	0x37, 0x43, 0x37, 0x08, 0x3D, 0x24, 0x43, 0x15, 0x5F, 0x05, 0x6D, 0x38,
	0x55, 0x25, 0x18, 0x36, 0x1C, 0x0F, 0x05, 0x1D, 0x05, 0x43, 0x39, 0x17,
	0x3D, 0x37, 0x39, 0x2E, 0x3A, 0x59, 0x14, 0x24, 0x14, 0x2D, 0x59, 0x32,
	0x1E, 0x2E, 0x24, 0x1F, 0x33, 0x0A, 0x10, 0x1E, 0x32, 0x6D, 0x5D, 0x52,
	0x23, 0x1D, 0x3B, 0x1D, 0x36, 0x36, 0x25, 0x28, 0x5B, 0x36, 0x20, 0x05,
	0x10, 0x1C, 0x0D, 0x18, 0x3E, 0x26, 0x02, 0x0F, 0x01, 0x3D, 0x73, 0x02,
	0x29, 0x36, 0x1F, 0x76, 0x0B, 0x04, 0x1E, 0x1A, 0x0A, 0x18, 0x11, 0x14,
	0x03, 0x31, 0x04, 0x04, 0x5E, 0x5B, 0x18, 0x07, 0x29, 0x06, 0x0A, 0x76,
	0x02, 0x08, 0x1E, 0x23, 0x38, 0x3C, 0x2A, 0x09, 0x13, 0x11, 0x09, 0x13,
	0x2D, 0x5F, 0x30, 0x54, 0x07, 0x58, 0x03, 0x75, 0x2A, 0x4E, 0x2F, 0x04,
	0x33, 0x1D, 0x33, 0x06, 0x0E, 0x06, 0x1D, 0x3B, 0x2D, 0x3A, 0x07, 0x3F,
	0x2E, 0x01, 0x2E, 0x07, 0x0B, 0x0F, 0x27, 0x31, 0x08, 0x3B, 0x06, 0x07,
	0x2A, 0x31, 0x01, 0x2A, 0x03, 0x03, 0x05, 0x3D, 0x25, 0x23, 0x13, 0x03,
	0x22, 0x51, 0x19, 0x0C, 0x23, 0x04, 0x33, 0x3B, 0x3D, 0x0A, 0x3F, 0x34,
	0x34, 0x39, 0x15, 0x3A, 0x09, 0x3F, 0x39, 0x18, 0x2A, 0x51, 0x20, 0x1C,
	0x18, 0x05, 0x32, 0x57, 0x3A, 0x35, 0x0A, 0x02, 0x16, 0x0F, 0x37, 0x19,
	0x14, 0x1C, 0x5D, 0x37, 0x5B, 0x13, 0x1F, 0x19, 0x27, 0x5F, 0x36, 0x36,
	0x5E, 0x23, 0x0E, 0x2C, 0x24, 0x24, 0x13, 0x2B, 0x20, 0x07, 0x2E, 0x0B,
	0x2E, 0x12, 0x27, 0x07, 0x1A, 0x23, 0x50, 0x21, 0x28, 0x0B, 0x25, 0x28,
	0x5B, 0x2F, 0x77, 0x0A, 0x37, 0x34, 0x58, 0x37, 0x19, 0x38, 0x3C, 0x2E,
	0x24, 0x0E, 0x4E, 0x00, 0x44, 0x6D, 0x43, 0x0F, 0x45, 0x0D, 0x17, 0x04,
	0x51, 0x5B, 0x0D, 0x16, 0x59, 0x50, 0x25, 0x05, 0x33, 0x07, 0x54, 0x38,
	0x05, 0x16, 0x1C, 0x37, 0x2D, 0x0E, 0x10, 0x3F, 0x17, 0x2D, 0x38, 0x00,
	0x15, 0x08, 0x58, 0x0C, 0x0B, 0x01, 0x59, 0x39, 0x5D, 0x17, 0x5B, 0x03,
	0x34, 0x1D, 0x20, 0x3F, 0x35, 0x2D, 0x40, 0x1A, 0x5C, 0x2C, 0x1B, 0x3B,
	0x73, 0x19, 0x17, 0x21, 0x53, 0x2A, 0x02, 0x12, 0x24, 0x3C, 0x37, 0x00,
	0x08, 0x26, 0x58, 0x08, 0x06, 0x06, 0x19, 0x18, 0x3B, 0x0D, 0x3B, 0x00,
	0x5D, 0x7B, 0x07, 0x29, 0x28, 0x52, 0x2B, 0x16, 0x39, 0x26, 0x19, 0x70,
	0x24, 0x17, 0x23, 0x5B, 0x18, 0x36, 0x57, 0x05, 0x38, 0x3A, 0x0E, 0x30,
	0x1D, 0x1C, 0x34, 0x21, 0x14, 0x5B, 0x3A, 0x77, 0x07, 0x17, 0x58, 0x2F,
	0x27, 0x36, 0x05, 0x1B, 0x53, 0x2A, 0x24, 0x04, 0x03, 0x06, 0x08, 0x19,
	0x54, 0x2B, 0x27, 0x2C, 0x3A, 0x36, 0x38, 0x3F, 0x0D, 0x58, 0x00, 0x28,
	0x53, 0x0C, 0x59, 0x4A, 0x58, 0x0C, 0x0A, 0x5E, 0x15, 0x27, 0x0C, 0x7B,
	0x3A, 0x36, 0x41, 0x0C, 0x13, 0x05, 0x04, 0x39, 0x31, 0x26, 0x23, 0x19,
	0x29, 0x52, 0x25, 0x29, 0x13, 0x57, 0x2A, 0x35, 0x19, 0x37, 0x04, 0x5C,
	0x24, 0x3A, 0x2C, 0x59, 0x5E, 0x34, 0x19, 0x04, 0x0A, 0x04, 0x7A, 0x14,
	0x0B, 0x5B, 0x3D, 0x0C, 0x28, 0x4A, 0x1B, 0x2A, 0x38, 0x38, 0x37, 0x01,
	0x22, 0x03, 0x07, 0x04, 0x03, 0x07, 0x75, 0x3F, 0x56, 0x3F, 0x11, 0x37,
	0x22, 0x14, 0x5E, 0x22, 0x26, 0x2B, 0x55, 0x29, 0x05, 0x70, 0x04, 0x26,
	0x01, 0x24, 0x0A, 0x36, 0x0D, 0x56, 0x0E, 0x25, 0x20, 0x4A, 0x07, 0x28,
	0x06, 0x3D, 0x52, 0x41, 0x3F, 0x0D, 0x1A, 0x29, 0x2C, 0x0F, 0x23, 0x3C,
	0x19, 0x59, 0x39, 0x20, 0x3C, 0x2F, 0x27, 0x21, 0x36, 0x43, 0x05, 0x1C,
	0x1F, 0x35, 0x02, 0x12, 0x0A, 0x1B, 0x18, 0x5E, 0x00, 0x5C, 0x0A, 0x71,
	0x3A, 0x14, 0x5E, 0x59, 0x25, 0x5B, 0x1B, 0x2A, 0x2F, 0x6D, 0x5A, 0x03,
	0x3F, 0x02, 0x30, 0x38, 0x33, 0x0F, 0x11, 0x69, 0x26, 0x24, 0x39, 0x44,
	0x11, 0x22, 0x2C, 0x18, 0x26, 0x09, 0x15, 0x18, 0x0D, 0x1E, 0x17, 0x04,
	0x07, 0x3F, 0x39, 0x0E, 0x55, 0x29, 0x03, 0x5C, 0x2D, 0x2E, 0x59, 0x20,
	0x1B, 0x33, 0x0D, 0x58, 0x05, 0x53, 0x34, 0x3F, 0x59, 0x3C, 0x2F, 0x0D,
	0x22, 0x06, 0x1F, 0x11, 0x16, 0x2F, 0x2F, 0x22, 0x22, 0x0F, 0x43, 0x16,
	0x28, 0x22, 0x26, 0x5F, 0x56, 0x2B, 0x0D, 0x71, 0x0F, 0x53, 0x16, 0x04,
	0x77, 0x1D, 0x08, 0x09, 0x1C, 0x6D, 0x5D, 0x00, 0x58, 0x0C, 0x15, 0x0A,
	0x14, 0x23, 0x28, 0x0F, 0x1E, 0x14, 0x3F, 0x1C, 0x3B, 0x21, 0x0C, 0x41,
	0x38, 0x31, 0x08, 0x23, 0x2D, 0x1F, 0x29, 0x35, 0x24, 0x0D, 0x12, 0x31,
	0x07, 0x33, 0x59, 0x19, 0x7B, 0x5E, 0x17, 0x0F, 0x09, 0x11, 0x5A, 0x56,
	0x22, 0x0F, 0x04, 0x19, 0x27, 0x59, 0x29, 0x20, 0x3F, 0x03, 0x1A, 0x0F,
	0x35, 0x01, 0x54, 0x0A, 0x59, 0x2F, 0x5C, 0x33, 0x1B, 0x44, 0x70, 0x00,
	0x05, 0x1C, 0x1E, 0x27, 0x5F, 0x33, 0x0F, 0x32, 0x05, 0x36, 0x51, 0x25,
	0x0F, 0x03, 0x38, 0x53, 0x2B, 0x13, 0x18, 0x1E, 0x26, 0x01, 0x26, 0x2A,
	0x0D, 0x2D, 0x56, 0x0D, 0x10, 0x3B, 0x0F, 0x14, 0x13, 0x76, 0x0D, 0x4E,
	0x22, 0x33, 0x15, 0x2A, 0x07, 0x18, 0x2E, 0x2F, 0x1B, 0x14, 0x26, 0x53,
	0x25, 0x47, 0x1B, 0x0D, 0x1C, 0x26, 0x07, 0x59, 0x22, 0x05, 0x25, 0x0F,
	0x3B, 0x09, 0x25, 0x73, 0x07, 0x53, 0x2D, 0x38, 0x05, 0x5A, 0x39, 0x2C,
	0x31, 0x0B, 0x29, 0x2E, 0x06, 0x28, 0x14, 0x3E, 0x0E, 0x0B, 0x3B, 0x24,
	0x47, 0x2E, 0x28, 0x05, 0x27, 0x3D, 0x32, 0x25, 0x1F, 0x26, 0x3D, 0x58,
	0x5B, 0x05, 0x74, 0x55, 0x06, 0x08, 0x04, 0x15, 0x54, 0x13, 0x1C, 0x3C,
	0x34, 0x07, 0x0B, 0x3F, 0x1D, 0x34, 0x04, 0x05, 0x26, 0x00, 0x24, 0x19,
	0x50, 0x0A, 0x19, 0x00, 0x2D, 0x0B, 0x23, 0x5D, 0x1B, 0x3F, 0x2E, 0x37,
	0x0A, 0x0D, 0x2A, 0x23, 0x59, 0x3B, 0x30, 0x18, 0x07, 0x17, 0x03, 0x04,
	0x1B, 0x14, 0x0F, 0x39, 0x70, 0x1C, 0x24, 0x0F, 0x0C, 0x76, 0x59, 0x00,
	0x39, 0x0C, 0x73, 0x5A, 0x38, 0x2F, 0x0C, 0x25, 0x35, 0x0C, 0x2F, 0x22,
	0x2F, 0x14, 0x29, 0x1E, 0x1F, 0x75, 0x28, 0x25, 0x3A, 0x59, 0x2E, 0x3D,
	0x27, 0x16, 0x59, 0x13, 0x2D, 0x59, 0x2F, 0x5F, 0x10, 0x5E, 0x11, 0x09,
	0x26, 0x3A, 0x27, 0x02, 0x5B, 0x06, 0x37, 0x5F, 0x57, 0x57, 0x05, 0x36,
	0x2D, 0x58, 0x1C, 0x1F, 0x27, 0x5C, 0x03, 0x07, 0x03, 0x14, 0x08, 0x17,
	0x34, 0x07, 0x00, 0x1F, 0x2C, 0x39, 0x22, 0x74, 0x3D, 0x36, 0x24, 0x39,
	0x10, 0x03, 0x50, 0x28, 0x18, 0x24, 0x25, 0x4E, 0x5E, 0x08, 0x30, 0x5B,
	0x53, 0x21, 0x58, 0x0C, 0x5E, 0x0C, 0x5E, 0x25, 0x37, 0x14, 0x53, 0x1B,
	0x58, 0x16, 0x0D, 0x16, 0x5C, 0x5B, 0x0A, 0x0D, 0x56, 0x3F, 0x3D, 0x70,
	0x5E, 0x50, 0x45, 0x5C, 0x0C, 0x36, 0x06, 0x37, 0x0F, 0x15, 0x1D, 0x52,
	0x2D, 0x0E, 0x35, 0x5E, 0x2C, 0x2B, 0x21, 0x06, 0x0D, 0x39, 0x0C, 0x09,
	0x0D, 0x03, 0x2A, 0x04, 0x0E, 0x1B, 0x1B, 0x50, 0x5E, 0x0A, 0x2C, 0x24,
	0x04, 0x5A, 0x32, 0x3A, 0x26, 0x22, 0x19, 0x59, 0x0F, 0x1A, 0x2A, 0x1C,
	0x26, 0x2A, 0x1E, 0x0E, 0x3E, 0x18, 0x1A, 0x29, 0x14, 0x1E, 0x0F, 0x2A,
	0x5C, 0x0C, 0x08, 0x3F, 0x33, 0x27, 0x27, 0x5D, 0x05, 0x1A, 0x5A, 0x09,
	0x29, 0x27, 0x14, 0x34, 0x00, 0x36, 0x1A, 0x18, 0x20, 0x2D, 0x06, 0x3A,
	0x0D, 0x19, 0x00, 0x17, 0x2C, 0x17, 0x47, 0x58, 0x2A, 0x59, 0x18, 0x54,
	0x06, 0x04, 0x5C, 0x28, 0x3E, 0x34, 0x34, 0x1F, 0x3A, 0x18, 0x02, 0x0C,
	0x1F, 0x10, 0x00, 0x29, 0x17, 0x2D, 0x11, 0x15, 0x55, 0x41, 0x5C, 0x12,
	0x5A, 0x09, 0x20, 0x2A, 0x29, 0x09, 0x28, 0x3A, 0x2C, 0x20, 0x0E, 0x56,
	0x04, 0x25, 0x33, 0x02, 0x2F, 0x0D, 0x0A, 0x35, 0x15, 0x36, 0x59, 0x3A,
	0x06, 0x1C, 0x23, 0x05, 0x0A, 0x08, 0x23, 0x58, 0x5B, 0x5A, 0x76, 0x19,
	0x54, 0x26, 0x21, 0x6D, 0x1B, 0x33, 0x04, 0x06, 0x21, 0x01, 0x59, 0x09,
	0x33, 0x71, 0x03, 0x09, 0x03, 0x12, 0x32, 0x20, 0x22, 0x26, 0x0E, 0x77,
	0x22, 0x55, 0x0B, 0x5C, 0x71, 0x23, 0x2C, 0x2F, 0x38, 0x27, 0x38, 0x30,
	0x25, 0x1B, 0x11, 0x1C, 0x16, 0x05, 0x02, 0x34, 0x47, 0x14, 0x2A, 0x03,
	0x04, 0x28, 0x57, 0x16, 0x3C, 0x0F, 0x43, 0x1B, 0x06, 0x27, 0x07, 0x20,
	0x0D, 0x20, 0x13, 0x12, 0x2D, 0x16, 0x2B, 0x1D, 0x2B, 0x5D, 0x4E, 0x09,
	0x00, 0x07, 0x58, 0x12, 0x5F, 0x22, 0x0F, 0x0F, 0x34, 0x3E, 0x1D, 0x18,
	0x23, 0x0B, 0x24, 0x39, 0x2E, 0x25, 0x2F, 0x25, 0x3E, 0x7A, 0x35, 0x56,
	0x59, 0x2A, 0x2B, 0x08, 0x09, 0x27, 0x1C, 0x33, 0x04, 0x24, 0x09, 0x39,
	0x3A, 0x5E, 0x20, 0x00, 0x44, 0x21, 0x5D, 0x28, 0x3B, 0x3A, 0x16, 0x1B,
	0x22, 0x38, 0x3A, 0x1B, 0x43, 0x09, 0x27, 0x3C, 0x76, 0x0F, 0x00, 0x5D,
	0x53, 0x16, 0x2F, 0x15, 0x21, 0x0A, 0x35, 0x21, 0x19, 0x1A, 0x2A, 0x38,
	0x5B, 0x00, 0x22, 0x23, 0x7B, 0x43, 0x1B, 0x2A, 0x38, 0x08, 0x55, 0x28,
	0x59, 0x2E, 0x72, 0x0B, 0x14, 0x0B, 0x33, 0x34, 0x3E, 0x0E, 0x21, 0x05,
	0x05, 0x3D, 0x59, 0x2F, 0x21, 0x34, 0x54, 0x54, 0x02, 0x31, 0x72, 0x29,
	0x0B, 0x3E, 0x0D, 0x26, 0x2D, 0x55, 0x23, 0x3F, 0x0D, 0x59, 0x27, 0x00,
	0x2F, 0x70, 0x22, 0x0E, 0x09, 0x2C, 0x15, 0x04, 0x0B, 0x05, 0x1A, 0x2D,
	0x2D, 0x51, 0x41, 0x32, 0x08, 0x3A, 0x07, 0x2F, 0x03, 0x27, 0x28, 0x02,
	0x07, 0x52, 0x26, 0x1E, 0x34, 0x59, 0x3B, 0x35, 0x1C, 0x07, 0x45, 0x2E,
	0x17, 0x0D, 0x0F, 0x59, 0x24, 0x7A, 0x34, 0x4E, 0x56, 0x01, 0x11, 0x16,
	0x0C, 0x28, 0x00, 0x0D, 0x59, 0x16, 0x29, 0x23, 0x71, 0x07, 0x12, 0x18,
	0x20, 0x69, 0x0D, 0x30, 0x0F, 0x02, 0x2F, 0x5C, 0x2E, 0x5F, 0x0D, 0x33,
	0x07, 0x22, 0x09, 0x18, 0x2A, 0x5C, 0x2C, 0x3D, 0x3C, 0x25, 0x3E, 0x2D,
	0x3A, 0x08, 0x07, 0x2A, 0x00, 0x39, 0x3D, 0x33, 0x1D, 0x08, 0x2A, 0x1F,
	0x2F, 0x3F, 0x50, 0x3E, 0x59, 0x2D, 0x55, 0x0F, 0x34, 0x0D, 0x7B, 0x2E,
	0x11, 0x21, 0x3D, 0x0B, 0x38, 0x30, 0x1B, 0x0E, 0x6D, 0x43, 0x3B, 0x21,
	0x2D, 0x04, 0x14, 0x0D, 0x1D, 0x3A, 0x09, 0x2B, 0x00, 0x34, 0x31, 0x23,
	0x00, 0x05, 0x0D, 0x24, 0x72, 0x36, 0x0D, 0x5F, 0x29, 0x72, 0x0D, 0x26,
	0x56, 0x38, 0x2C, 0x1E, 0x15, 0x06, 0x26, 0x3B, 0x0A, 0x34, 0x2D, 0x0D,
	0x7A, 0x35, 0x0A, 0x22, 0x27, 0x38, 0x0B, 0x12, 0x59, 0x3A, 0x15, 0x5B,
	0x17, 0x38, 0x02, 0x2E, 0x2A, 0x4A, 0x1C, 0x22, 0x00, 0x3C, 0x24, 0x03,
	0x44, 0x28, 0x5B, 0x0E, 0x23, 0x03, 0x70, 0x25, 0x52, 0x5A, 0x21, 0x10,
	0x0D, 0x10, 0x3A, 0x21, 0x27, 0x29, 0x4A, 0x26, 0x5C, 0x23, 0x0D, 0x19,
	0x05, 0x44, 0x00, 0x2E, 0x22, 0x23, 0x21, 0x73, 0x00, 0x0F, 0x34, 0x52,
	0x11, 0x0A, 0x09, 0x37, 0x2C, 0x2C, 0x1A, 0x35, 0x5C, 0x1C, 0x11, 0x15,
	0x32, 0x1E, 0x26, 0x08, 0x20, 0x0D, 0x2F, 0x00, 0x33, 0x16, 0x35, 0x5F,
	0x0D, 0x77, 0x19, 0x2B, 0x2F, 0x21, 0x15, 0x01, 0x04, 0x21, 0x5B, 0x33,
	0x07, 0x25, 0x19, 0x0E, 0x03, 0x25, 0x0D, 0x2C, 0x28, 0x14, 0x25, 0x16,
	0x17, 0x18, 0x70, 0x3A, 0x2E, 0x00, 0x31, 0x01, 0x3C, 0x12, 0x23, 0x03,
	0x2C, 0x0F, 0x30, 0x21, 0x05, 0x34, 0x47, 0x02, 0x27, 0x1B, 0x6D, 0x54,
	0x56, 0x36, 0x19, 0x0D, 0x29, 0x22, 0x5A, 0x21, 0x03, 0x24, 0x0D, 0x1D,
	0x5B, 0x2A, 0x0D, 0x53, 0x08, 0x5C, 0x00, 0x5D, 0x54, 0x5F, 0x3E, 0x2D,
	0x25, 0x36, 0x14, 0x2D, 0x0D, 0x2D, 0x38, 0x39, 0x5C, 0x0F, 0x1A, 0x0F,
	0x04, 0x53, 0x12, 0x0A, 0x2B, 0x14, 0x39, 0x2A, 0x1B, 0x59, 0x0B, 0x20,
	0x0E, 0x20, 0x14, 0x0B, 0x32, 0x77, 0x55, 0x36, 0x58, 0x0A, 0x36, 0x21,
	0x0F, 0x38, 0x31, 0x0A, 0x28, 0x02, 0x0B, 0x32, 0x20, 0x1B, 0x2E, 0x45,
	0x04, 0x09, 0x02, 0x23, 0x29, 0x3B, 0x6D, 0x27, 0x10, 0x5D, 0x06, 0x00,
	0x1B, 0x2E, 0x37, 0x2E, 0x1A, 0x0A, 0x33, 0x09, 0x22, 0x05, 0x25, 0x13,
	0x18, 0x5F, 0x7A, 0x20, 0x24, 0x17, 0x29, 0x33, 0x19, 0x25, 0x2D, 0x29,
	0x2D, 0x35, 0x29, 0x0A, 0x31, 0x07, 0x2E, 0x56, 0x1D, 0x0F, 0x24, 0x38,
	0x02, 0x0D, 0x18, 0x3A, 0x1A, 0x57, 0x3E, 0x01, 0x2E, 0x05, 0x15, 0x1E,
	0x3E, 0x16, 0x09, 0x2F, 0x06, 0x01, 0x36, 0x00, 0x19, 0x3A, 0x52, 0x35,
	0x3A, 0x28, 0x59, 0x3E, 0x00, 0x35, 0x22, 0x5D, 0x20, 0x20, 0x43, 0x35,
	0x1E, 0x0A, 0x0B, 0x39, 0x30, 0x38, 0x04, 0x11, 0x1D, 0x59, 0x14, 0x44,
	0x04, 0x25, 0x31, 0x09, 0x5E, 0x15, 0x23, 0x16, 0x04, 0x1D, 0x29, 0x35,
	0x04, 0x09, 0x26, 0x76, 0x1F, 0x55, 0x2B, 0x04, 0x69, 0x38, 0x51, 0x29,
	0x3C, 0x25, 0x3C, 0x2C, 0x3A, 0x01, 0x75, 0x2F, 0x4A, 0x07, 0x3B, 0x36,
	0x34, 0x13, 0x03, 0x2D, 0x17, 0x3D, 0x0C, 0x03, 0x23, 0x2A, 0x23, 0x02,
	0x39, 0x03, 0x76, 0x5D, 0x2D, 0x0F, 0x40, 0x18, 0x1C, 0x54, 0x37, 0x1D,
	0x27, 0x36, 0x0F, 0x2A, 0x5C, 0x0C, 0x47, 0x02, 0x1F, 0x5F, 0x71, 0x06,
	0x52, 0x0C, 0x0F, 0x07, 0x39, 0x37, 0x39, 0x09, 0x7B, 0x27, 0x10, 0x23,
	0x58, 0x0D, 0x35, 0x51, 0x0C, 0x0E, 0x32, 0x54, 0x53, 0x04, 0x3B, 0x00,
	0x5F, 0x53, 0x2C, 0x59, 0x7B, 0x3C, 0x34, 0x3C, 0x0A, 0x0E, 0x24, 0x53,
	0x39, 0x44, 0x69, 0x03, 0x0F, 0x3F, 0x2F, 0x14, 0x58, 0x02, 0x2C, 0x22,
	0x2E, 0x54, 0x26, 0x2C, 0x03, 0x17, 0x5F, 0x2B, 0x24, 0x09, 0x2C, 0x2D,
	0x27, 0x37, 0x01, 0x2B, 0x3C, 0x39, 0x45, 0x2F, 0x3A, 0x1E, 0x19, 0x24,
	0x1F, 0x71, 0x02, 0x56, 0x38, 0x59, 0x23, 0x02, 0x2C, 0x25, 0x3F, 0x03,
	0x1A, 0x32, 0x0F, 0x18, 0x7B, 0x0D, 0x33, 0x34, 0x1B, 0x77, 0x5C, 0x16,
	0x3E, 0x29, 0x0A, 0x5A, 0x56, 0x07, 0x3A, 0x03, 0x58, 0x59, 0x28, 0x59,
	0x32, 0x0A, 0x33, 0x2A, 0x03, 0x07, 0x1E, 0x59, 0x16, 0x21, 0x15, 0x29,
	0x0A, 0x16, 0x1F, 0x72, 0x5E, 0x0C, 0x02, 0x44, 0x01, 0x5C, 0x4E, 0x23,
	0x21, 0x2B, 0x05, 0x52, 0x41, 0x27, 0x29, 0x20, 0x34, 0x0B, 0x23, 0x3B,
	0x39, 0x2B, 0x1C, 0x2D, 0x3B, 0x3B, 0x17, 0x16, 0x08, 0x10, 0x03, 0x56,
	0x19, 0x0C, 0x69, 0x00, 0x22, 0x1A, 0x5F, 0x2B, 0x2F, 0x33, 0x01, 0x01,
	0x26, 0x2B, 0x27, 0x1B, 0x0A, 0x0A, 0x0D, 0x06, 0x3E, 0x5F, 0x72, 0x08,
	0x57, 0x27, 0x0D, 0x1A, 0x15, 0x4A, 0x2B, 0x5A, 0x32, 0x35, 0x0B, 0x29,
	0x08, 0x6D, 0x5C, 0x16, 0x29, 0x11, 0x24, 0x22, 0x54, 0x02, 0x02, 0x2F,
	0x0D, 0x29, 0x0F, 0x53, 0x12, 0x5C, 0x51, 0x41, 0x58, 0x32, 0x43, 0x26,
	0x04, 0x1D, 0x24, 0x28, 0x27, 0x19, 0x5E, 0x15, 0x58, 0x34, 0x0A, 0x2F,
	0x33, 0x3F, 0x20, 0x59, 0x5C, 0x03, 0x47, 0x31, 0x06, 0x5C, 0x0D, 0x27,
	0x53, 0x24, 0x07, 0x6D, 0x1D, 0x2E, 0x06, 0x26, 0x06, 0x1E, 0x50, 0x00,
	0x39, 0x6D, 0x43, 0x09, 0x18, 0x3A, 0x29, 0x43, 0x36, 0x59, 0x5B, 0x06,
	0x3D, 0x16, 0x5B, 0x2E, 0x18, 0x26, 0x54, 0x03, 0x2A, 0x23, 0x3A, 0x12,
	0x23, 0x20, 0x16, 0x22, 0x0C, 0x3E, 0x1A, 0x1A, 0x3D, 0x17, 0x25, 0x5A,
	0x32, 0x02, 0x22, 0x37, 0x52, 0x2C, 0x0E, 0x2B, 0x20, 0x2C, 0x72, 0x18,
	0x0C, 0x2B, 0x31, 0x2D, 0x2B, 0x0B, 0x1B, 0x3E, 0x0E, 0x3F, 0x0B, 0x14,
	0x1B, 0x2E, 0x29, 0x25, 0x45, 0x0F, 0x03, 0x2D, 0x30, 0x2F, 0x12, 0x32,
	0x06, 0x00, 0x39, 0x05, 0x00, 0x59, 0x56, 0x21, 0x0C, 0x0E, 0x04, 0x28,
	0x0B, 0x5F, 0x13, 0x35, 0x18, 0x5E, 0x2A, 0x09, 0x34, 0x54, 0x56, 0x0F,
	0x3A, 0x2D, 0x34, 0x24, 0x28, 0x04, 0x55, 0x12, 0x3D, 0x28, 0x71, 0x3B,
	0x10, 0x07, 0x52, 0x01, 0x28, 0x55, 0x28, 0x23, 0x24, 0x5E, 0x38, 0x19,
	0x3E, 0x0C, 0x36, 0x26, 0x27, 0x24, 0x7A, 0x21, 0x19, 0x08, 0x2A, 0x69,
	0x0A, 0x09, 0x21, 0x0D, 0x2F, 0x3D, 0x35, 0x3B, 0x0F, 0x11, 0x08, 0x2E,
	0x57, 0x1F, 0x75, 0x5F, 0x15, 0x2F, 0x2A, 0x0F, 0x05, 0x17, 0x17, 0x07,
	0x0A, 0x0B, 0x30, 0x1C, 0x18, 0x31, 0x43, 0x53, 0x02, 0x2C, 0x37, 0x5A,
	0x0E, 0x41, 0x3E, 0x75, 0x22, 0x18, 0x39, 0x02, 0x71, 0x55, 0x12, 0x0D,
	0x3D, 0x04, 0x2F, 0x38, 0x1E, 0x0C, 0x15, 0x47, 0x14, 0x1C, 0x09, 0x24,
	0x2B, 0x27, 0x20, 0x27, 0x27, 0x14, 0x12, 0x0F, 0x0C, 0x32, 0x03, 0x37,
	0x29, 0x08, 0x00, 0x04, 0x17, 0x0B, 0x2A, 0x74, 0x00, 0x51, 0x37, 0x5E,
	0x10, 0x0D, 0x26, 0x04, 0x2C, 0x26, 0x2F, 0x24, 0x23, 0x1E, 0x36, 0x43,
	0x55, 0x29, 0x06, 0x2D, 0x0B, 0x29, 0x38, 0x1E, 0x09, 0x20, 0x32, 0x2A,
	0x18, 0x12, 0x1E, 0x02, 0x24, 0x07, 0x2D, 0x43, 0x26, 0x24, 0x31, 0x74,
	0x1E, 0x02, 0x2A, 0x12, 0x26, 0x01, 0x29, 0x19, 0x07, 0x0B, 0x23, 0x14,
	0x2B, 0x12, 0x0C, 0x59, 0x2F, 0x58, 0x5F, 0x28, 0x39, 0x10, 0x02, 0x3D,
	0x7A, 0x07, 0x17, 0x02, 0x07, 0x09, 0x1E, 0x23, 0x5D, 0x58, 0x2B, 0x55,
	0x57, 0x17, 0x39, 0x34, 0x07, 0x57, 0x0A, 0x2C, 0x1B, 0x3B, 0x20, 0x3F,
	0x06, 0x07, 0x36, 0x03, 0x25, 0x09, 0x38, 0x5E, 0x10, 0x5A, 0x05, 0x69,
	0x14, 0x13, 0x5B, 0x59, 0x23, 0x35, 0x4A, 0x38, 0x5E, 0x17, 0x5D, 0x16,
	0x00, 0x3D, 0x38, 0x00, 0x03, 0x5A, 0x5E, 0x26, 0x05, 0x31, 0x03, 0x0C,
	0x2D, 0x00, 0x50, 0x00, 0x0C, 0x0B, 0x59, 0x36, 0x56, 0x0D, 0x1B, 0x5E,
	0x0B, 0x23, 0x23, 0x70, 0x29, 0x4A, 0x3F, 0x3C, 0x2E, 0x2D, 0x51, 0x38,
	0x39, 0x17, 0x54, 0x2C, 0x38, 0x5F, 0x09, 0x3A, 0x36, 0x1F, 0x3E, 0x26,
	0x2A, 0x03, 0x0C, 0x3E, 0x69, 0x3E, 0x0F, 0x39, 0x5C, 0x16, 0x0B, 0x16,
	0x0B, 0x59, 0x23, 0x16, 0x05, 0x08, 0x3D, 0x32, 0x26, 0x24, 0x02, 0x33,
	0x23, 0x1B, 0x2D, 0x18, 0x05, 0x31, 0x16, 0x09, 0x3C, 0x38, 0x09, 0x43,
	0x54, 0x06, 0x03, 0x3B, 0x24, 0x29, 0x00, 0x5F, 0x71, 0x05, 0x26, 0x0D,
	0x1C, 0x11, 0x1E, 0x15, 0x00, 0x24, 0x0C, 0x21, 0x4A, 0x05, 0x5B, 0x0D,
	0x08, 0x58, 0x09, 0x0A, 0x0D, 0x20, 0x0D, 0x19, 0x1D, 0x23, 0x1F, 0x50,
	0x06, 0x05, 0x26, 0x43, 0x06, 0x14, 0x1A, 0x3A, 0x55, 0x4A, 0x2B, 0x3E,
	0x2B, 0x03, 0x52, 0x5B, 0x39, 0x09, 0x16, 0x04, 0x14, 0x00, 0x24, 0x1B,
	0x4A, 0x2A, 0x24, 0x01, 0x1C, 0x0B, 0x14, 0x5E, 0x06, 0x1A, 0x09, 0x3B,
	0x53, 0x0C, 0x38, 0x1B, 0x26, 0x07, 0x26, 0x0A, 0x26, 0x21, 0x05, 0x72,
	0x26, 0x2E, 0x45, 0x01, 0x09, 0x36, 0x18, 0x2D, 0x2A, 0x13, 0x2B, 0x35,
	0x3B, 0x5A, 0x2E, 0x2D, 0x16, 0x3E, 0x44, 0x03, 0x20, 0x1B, 0x41, 0x12,
	0x70, 0x02, 0x08, 0x2F, 0x2F, 0x75, 0x54, 0x07, 0x26, 0x0C, 0x69, 0x3D,
	0x05, 0x57, 0x40, 0x20, 0x05, 0x08, 0x1A, 0x24, 0x09, 0x2F, 0x03, 0x09,
	0x1A, 0x12, 0x5E, 0x26, 0x00, 0x06, 0x0B, 0x2F, 0x37, 0x18, 0x27, 0x37,
	0x34, 0x00, 0x23, 0x26, 0x2D, 0x36, 0x08, 0x2F, 0x5E, 0x23, 0x2B, 0x38,
	0x09, 0x2C, 0x72, 0x35, 0x24, 0x41, 0x29, 0x21, 0x20, 0x34, 0x14, 0x07,
	0x21, 0x5C, 0x0D, 0x27, 0x2C, 0x25, 0x04, 0x56, 0x01, 0x2A, 0x05, 0x0F,
	0x08, 0x09, 0x0C, 0x23, 0x03, 0x31, 0x09, 0x0F, 0x20, 0x2F, 0x33, 0x59,
	0x2F, 0x0D, 0x29, 0x30, 0x25, 0x52, 0x15, 0x2D, 0x3B, 0x1C, 0x31, 0x2C,
	0x2E, 0x10, 0x14, 0x40, 0x10, 0x1C, 0x2C, 0x29, 0x26, 0x37, 0x1A, 0x37,
	0x39, 0x1A, 0x34, 0x1E, 0x2B, 0x29, 0x0E, 0x1A, 0x28, 0x08, 0x2A, 0x1C,
	0x12, 0x2B, 0x34, 0x3B, 0x27, 0x27, 0x3B, 0x3B, 0x28, 0x24, 0x7A, 0x1A,
	0x1B, 0x3C, 0x01, 0x0C, 0x16, 0x2F, 0x5E, 0x3B, 0x26, 0x28, 0x24, 0x1A,
	0x2C, 0x36, 0x1C, 0x39, 0x26, 0x5A, 0x08, 0x1F, 0x26, 0x5E, 0x40, 0x03,
	0x20, 0x56, 0x00, 0x1B, 0x0E, 0x02, 0x06, 0x58, 0x22, 0x3B, 0x2F, 0x50,
	0x1B, 0x07, 0x32, 0x05, 0x0D, 0x07, 0x0F, 0x10, 0x29, 0x0D, 0x14, 0x1B,
	0x31, 0x2F, 0x2E, 0x57, 0x3D, 0x0A, 0x2F, 0x50, 0x2A, 0x0E, 0x06, 0x34,
	0x31, 0x27, 0x2F, 0x3B, 0x00, 0x4E, 0x3E, 0x19, 0x38, 0x22, 0x11, 0x09,
	0x3B, 0x0A, 0x18, 0x4A, 0x01, 0x12, 0x71, 0x36, 0x38, 0x24, 0x24, 0x38,
	0x0A, 0x18, 0x56, 0x27, 0x06, 0x08, 0x00, 0x07, 0x07, 0x37, 0x1A, 0x55,
	0x1F, 0x0D, 0x77, 0x05, 0x28, 0x17, 0x31, 0x0C, 0x58, 0x33, 0x17, 0x3C,
	0x29, 0x1B, 0x34, 0x00, 0x1B, 0x2E, 0x35, 0x38, 0x3C, 0x59, 0x2E, 0x55,
	0x4E, 0x06, 0x39, 0x17, 0x22, 0x13, 0x39, 0x0F, 0x0F, 0x03, 0x13, 0x0C,
	0x26, 0x04, 0x3F, 0x2A, 0x27, 0x11, 0x14, 0x34, 0x29, 0x37, 0x2A, 0x00,
	0x3A, 0x12, 0x3E, 0x1E, 0x0F, 0x1B, 0x2D, 0x58, 0x1D, 0x10, 0x5D, 0x0B,
	0x0D, 0x5F, 0x75, 0x24, 0x05, 0x23, 0x1A, 0x03, 0x21, 0x2B, 0x58, 0x09,
	0x7A, 0x27, 0x2B, 0x5F, 0x22, 0x0E, 0x43, 0x0C, 0x1C, 0x5E, 0x2B, 0x01,
	0x36, 0x2B, 0x5F, 0x27, 0x21, 0x33, 0x06, 0x22, 0x34, 0x5D, 0x11, 0x19,
	0x2C, 0x2C, 0x54, 0x0D, 0x0D, 0x2F, 0x15, 0x2E, 0x23, 0x01, 0x1B, 0x38,
	0x47, 0x2C, 0x1D, 0x3E, 0x14, 0x5E, 0x12, 0x08, 0x58, 0x2C, 0x5D, 0x03,
	0x02, 0x2E, 0x05, 0x20, 0x17, 0x16, 0x1E, 0x2E, 0x3D, 0x4A, 0x1D, 0x2E,
	0x16, 0x0A, 0x0F, 0x19, 0x0A, 0x21, 0x01, 0x02, 0x20, 0x1D, 0x70, 0x09,
	0x30, 0x3E, 0x5E, 0x0B, 0x3D, 0x04, 0x08, 0x02, 0x10, 0x38, 0x06, 0x5B,
	0x23, 0x32, 0x3A, 0x2E, 0x58, 0x2A, 0x69, 0x43, 0x20, 0x0D, 0x1D, 0x25,
	0x54, 0x37, 0x5F, 0x2E, 0x2B, 0x39, 0x2B, 0x2B, 0x02, 0x10, 0x0D, 0x4A,
	0x34, 0x25, 0x7B, 0x03, 0x08, 0x00, 0x52, 0x15, 0x21, 0x17, 0x06, 0x06,
	0x2F, 0x27, 0x2E, 0x2F, 0x1B, 0x17, 0x34, 0x25, 0x06, 0x5D, 0x7A, 0x26,
	0x29, 0x5C, 0x0A, 0x7B, 0x2A, 0x55, 0x05, 0x3B, 0x26, 0x55, 0x16, 0x3B,
	0x02, 0x13, 0x47, 0x25, 0x57, 0x07, 0x70, 0x28, 0x25, 0x5A, 0x3E, 0x32,
	0x2B, 0x2B, 0x18, 0x3D, 0x34, 0x0A, 0x36, 0x29, 0x05, 0x34, 0x24, 0x09,
	0x23, 0x24, 0x0E, 0x28, 0x24, 0x38, 0x29, 0x36, 0x27, 0x33, 0x07, 0x12,
	0x04, 0x02, 0x07, 0x37, 0x5A, 0x10, 0x1E, 0x2F, 0x1B, 0x53, 0x26, 0x06,
	0x30, 0x00, 0x0F, 0x69, 0x47, 0x18, 0x56, 0x31, 0x1B, 0x06, 0x4A, 0x01,
	0x2E, 0x77, 0x2E, 0x56, 0x2D, 0x23, 0x18, 0x09, 0x00, 0x06, 0x3C, 0x2E,
	0x3A, 0x0A, 0x26, 0x20, 0x16, 0x54, 0x53, 0x19, 0x32, 0x24, 0x03, 0x34,
	0x5A, 0x0E, 0x2D, 0x04, 0x0C, 0x59, 0x3A, 0x1B, 0x2E, 0x2B, 0x03, 0x25,
	0x27, 0x0D, 0x0F, 0x14, 0x13, 0x23, 0x1A, 0x56, 0x1D, 0x04, 0x31, 0x14,
	0x14, 0x2D, 0x22, 0x34, 0x5B, 0x23, 0x36, 0x52, 0x74, 0x04, 0x35, 0x02,
	0x3B, 0x75, 0x47, 0x20, 0x58, 0x1F, 0x26, 0x2E, 0x58, 0x34, 0x0C, 0x2F,
	0x5E, 0x37, 0x5E, 0x21, 0x6D, 0x25, 0x0F, 0x41, 0x5C, 0x7A, 0x21, 0x11,
	0x58, 0x1A, 0x76, 0x23, 0x29, 0x08, 0x5D, 0x01, 0x55, 0x56, 0x5A, 0x3E,
	0x74, 0x15, 0x3B, 0x03, 0x28, 0x1A, 0x27, 0x0A, 0x22, 0x07, 0x0A, 0x15,
	0x0D, 0x59, 0x2A, 0x1B, 0x23, 0x08, 0x1D, 0x1C, 0x21, 0x3C, 0x0E, 0x3D,
	0x28, 0x2D, 0x16, 0x04, 0x24, 0x27, 0x15, 0x26, 0x4E, 0x06, 0x0A, 0x38,
	0x34, 0x00, 0x1F, 0x00, 0x74, 0x24, 0x08, 0x5F, 0x3A, 0x71, 0x3A, 0x55,
	0x01, 0x58, 0x17, 0x2F, 0x55, 0x56, 0x3C, 0x0C, 0x3E, 0x36, 0x5C, 0x44,
	0x77, 0x2B, 0x38, 0x25, 0x1E, 0x2E, 0x06, 0x31, 0x1B, 0x5B, 0x24, 0x5C,
	0x38, 0x39, 0x29, 0x7B, 0x20, 0x0E, 0x38, 0x19, 0x31, 0x3F, 0x08, 0x19,
	0x18, 0x31, 0x20, 0x55, 0x3B, 0x3C, 0x23, 0x5B, 0x32, 0x20, 0x1E, 0x16,
	0x2B, 0x0B, 0x5B, 0x13, 0x38, 0x3E, 0x3B, 0x28, 0x0C, 0x69, 0x54, 0x3B,
	0x09, 0x06, 0x6D, 0x38, 0x14, 0x5B, 0x23, 0x35, 0x16, 0x04, 0x16, 0x2C,
	0x20, 0x59, 0x4E, 0x1B, 0x1D, 0x13, 0x0D, 0x4A, 0x14, 0x11, 0x0A, 0x58,
	0x17, 0x00, 0x0A, 0x16, 0x03, 0x02, 0x0D, 0x32, 0x2C, 0x2D, 0x35, 0x08,
	0x07, 0x24, 0x2D, 0x3B, 0x38, 0x5E, 0x2B, 0x07, 0x32, 0x03, 0x03, 0x0B,
	0x03, 0x25, 0x06, 0x58, 0x06, 0x27, 0x13, 0x1B, 0x1D, 0x75, 0x2F, 0x55,
	0x1C, 0x2D, 0x18, 0x34, 0x32, 0x14, 0x38, 0x0E, 0x20, 0x28, 0x00, 0x2F,
	0x00, 0x55, 0x56, 0x03, 0x2A, 0x74, 0x16, 0x09, 0x1E, 0x0A, 0x21, 0x2D,
	0x51, 0x00, 0x32, 0x71, 0x06, 0x26, 0x5E, 0x40, 0x25, 0x1A, 0x1B, 0x1F,
	0x08, 0x23, 0x2E, 0x04, 0x24, 0x33, 0x72, 0x14, 0x58, 0x00, 0x29, 0x69,
	0x5A, 0x06, 0x01, 0x23, 0x35, 0x2B, 0x04, 0x24, 0x0F, 0x0C, 0x3D, 0x09,
	0x2C, 0x3F, 0x06, 0x25, 0x2A, 0x3F, 0x23, 0x2E, 0x1F, 0x54, 0x28, 0x32,
	0x25, 0x14, 0x57, 0x56, 0x53, 0x15, 0x25, 0x27, 0x05, 0x12, 0x6D, 0x2B,
	0x2A, 0x1F, 0x0A, 0x6D, 0x2D, 0x2E, 0x09, 0x33, 0x25, 0x43, 0x25, 0x20,
	0x22, 0x12, 0x36, 0x02, 0x2D, 0x04, 0x0A, 0x2F, 0x4E, 0x3B, 0x08, 0x06,
	0x2D, 0x59, 0x03, 0x5C, 0x06, 0x29, 0x15, 0x06, 0x2F, 0x03, 0x1B, 0x37,
	0x0C, 0x0F, 0x74, 0x2A, 0x06, 0x27, 0x18, 0x70, 0x3F, 0x16, 0x20, 0x0D,
	0x31, 0x06, 0x52, 0x38, 0x3A, 0x0C, 0x29, 0x28, 0x3D, 0x44, 0x30, 0x05,
	0x13, 0x1B, 0x31, 0x74, 0x23, 0x52, 0x0D, 0x0A, 0x0A, 0x1D, 0x58, 0x1F,
	0x2A, 0x1B, 0x06, 0x0D, 0x21, 0x26, 0x7A, 0x2E, 0x19, 0x26, 0x32, 0x30,
	0x01, 0x58, 0x45, 0x21, 0x2A, 0x22, 0x08, 0x03, 0x09, 0x2A, 0x2E, 0x03,
	0x18, 0x0A, 0x21, 0x5B, 0x19, 0x29, 0x11, 0x11, 0x3D, 0x06, 0x2C, 0x31,
	0x01, 0x47, 0x59, 0x45, 0x07, 0x12, 0x58, 0x58, 0x22, 0x2E, 0x30, 0x0F,
	0x30, 0x17, 0x12, 0x09, 0x58, 0x02, 0x08, 0x1A, 0x26, 0x0B, 0x19, 0x0A,
	0x13, 0x0A, 0x18, 0x0C, 0x2C, 0x32, 0x12, 0x3A, 0x18, 0x59, 0x0D, 0x0A,
	0x14, 0x0F, 0x21, 0x2C, 0x30, 0x3F, 0x1B, 0x03, 0x5B, 0x0B, 0x02, 0x52,
	0x5E, 0x3F, 0x10, 0x3B, 0x14, 0x36, 0x29, 0x7B, 0x18, 0x56, 0x04, 0x5F,
	0x37, 0x5F, 0x02, 0x0C, 0x1C, 0x37, 0x3C, 0x08, 0x1F, 0x58, 0x0A, 0x18,
	0x36, 0x1E, 0x1C, 0x28, 0x3A, 0x59, 0x1D, 0x2A, 0x6D, 0x1C, 0x36, 0x56,
	0x00, 0x18, 0x0B, 0x0F, 0x29, 0x20, 0x11, 0x34, 0x12, 0x3F, 0x0D, 0x31,
	0x24, 0x2A, 0x17, 0x0D, 0x05, 0x27, 0x0B, 0x3E, 0x58, 0x70, 0x05, 0x24,
	0x2C, 0x5D, 0x0D, 0x43, 0x15, 0x22, 0x25, 0x35, 0x21, 0x34, 0x08, 0x18,
	0x05, 0x27, 0x07, 0x5A, 0x1B, 0x12, 0x29, 0x32, 0x41, 0x58, 0x3B, 0x09,
	0x22, 0x34, 0x40, 0x17, 0x1B, 0x13, 0x45, 0x0F, 0x01, 0x43, 0x0C, 0x21,
	0x08, 0x34, 0x05, 0x52, 0x0F, 0x12, 0x04, 0x0A, 0x15, 0x5C, 0x26, 0x2A,
	0x02, 0x50, 0x45, 0x13, 0x29, 0x27, 0x4A, 0x18, 0x3C, 0x31, 0x0B, 0x07,
	0x06, 0x58, 0x26, 0x22, 0x07, 0x04, 0x5C, 0x10, 0x05, 0x2D, 0x02, 0x39,
	0x07, 0x00, 0x25, 0x0D, 0x19, 0x77, 0x36, 0x00, 0x36, 0x2A, 0x72, 0x34,
	0x11, 0x28, 0x21, 0x29, 0x14, 0x4E, 0x56, 0x0A, 0x10, 0x0E, 0x0A, 0x08,
	0x44, 0x16, 0x0E, 0x3B, 0x29, 0x19, 0x03, 0x05, 0x15, 0x59, 0x1D, 0x34,
	0x29, 0x0D, 0x57, 0x04, 0x2F, 0x01, 0x4E, 0x26, 0x3C, 0x09, 0x3F, 0x27,
	0x0B, 0x08, 0x2C, 0x58, 0x05, 0x41, 0x02, 0x28, 0x5B, 0x22, 0x5B, 0x40,
	0x0B, 0x0E, 0x39, 0x0B, 0x2A, 0x24, 0x3A, 0x50, 0x3F, 0x2D, 0x36, 0x5D,
	0x3B, 0x0A, 0x28, 0x3A, 0x09, 0x0C, 0x07, 0x05, 0x0E, 0x20, 0x16, 0x0A,
	0x00, 0x09, 0x1D, 0x2C, 0x09, 0x5D, 0x11, 0x08, 0x13, 0x1E, 0x26, 0x36,
	0x34, 0x28, 0x5D, 0x19, 0x00, 0x24, 0x22, 0x07, 0x08, 0x3B, 0x3E, 0x33,
	0x38, 0x0C, 0x07, 0x2E, 0x19, 0x09, 0x24, 0x0A, 0x02, 0x31, 0x02, 0x5C,
	0x15, 0x2F, 0x0C, 0x2C, 0x39, 0x20, 0x36, 0x04, 0x34, 0x40, 0x15, 0x02,
	0x50, 0x06, 0x3A, 0x2C, 0x55, 0x3B, 0x0A, 0x11, 0x0D, 0x39, 0x12, 0x0C,
	0x27, 0x73, 0x08, 0x30, 0x1F, 0x3D, 0x32, 0x47, 0x0E, 0x19, 0x3B, 0x77,
	0x1D, 0x20, 0x07, 0x07, 0x30, 0x24, 0x10, 0x1E, 0x1A, 0x37, 0x27, 0x55,
	0x3F, 0x33, 0x08, 0x19, 0x27, 0x24, 0x31, 0x74, 0x5B, 0x55, 0x0A, 0x20,
	0x10, 0x3A, 0x17, 0x0F, 0x33, 0x2B, 0x1E, 0x59, 0x5D, 0x03, 0x08, 0x2B,
	0x18, 0x5F, 0x0E, 0x04, 0x54, 0x56, 0x45, 0x58, 0x2A, 0x2D, 0x0F, 0x1F,
	0x1E, 0x09, 0x19, 0x52, 0x2B, 0x02, 0x77, 0x0A, 0x25, 0x2C, 0x38, 0x3B,
	0x18, 0x2D, 0x17, 0x3E, 0x0B, 0x1E, 0x16, 0x24, 0x3A, 0x38, 0x26, 0x23,
	0x09, 0x0A, 0x2F, 0x43, 0x0D, 0x5C, 0x0F, 0x33, 0x38, 0x29, 0x57, 0x0D,
	0x21, 0x3A, 0x28, 0x5E, 0x08, 0x07, 0x3E, 0x08, 0x57, 0x5B, 0x16, 0x1F,
	0x03, 0x5F, 0x12, 0x2C, 0x0F, 0x55, 0x21, 0x1F, 0x00, 0x1F, 0x38, 0x57,
	0x09, 0x70, 0x0B, 0x27, 0x21, 0x3F, 0x37, 0x21, 0x4E, 0x20, 0x24, 0x0A,
	0x21, 0x50, 0x16, 0x0D, 0x2A, 0x22, 0x54, 0x5B, 0x5F, 0x71, 0x1D, 0x06,
	0x41, 0x59, 0x20, 0x2F, 0x54, 0x1F, 0x09, 0x24, 0x3E, 0x0C, 0x24, 0x11,
	0x6D, 0x3C, 0x23, 0x1B, 0x52, 0x0E, 0x47, 0x13, 0x20, 0x44, 0x33, 0x0A,
	0x00, 0x23, 0x0A, 0x11, 0x21, 0x38, 0x04, 0x26, 0x13, 0x3C, 0x30, 0x37,
	0x52, 0x08, 0x05, 0x08, 0x5F, 0x0C, 0x0B, 0x01, 0x13, 0x57, 0x19, 0x04,
	0x05, 0x2D, 0x45, 0x00, 0x08, 0x0F, 0x09, 0x08, 0x26, 0x1A, 0x26, 0x11,
	0x2C, 0x1F, 0x2F, 0x39, 0x09, 0x06, 0x44, 0x32, 0x16, 0x53, 0x02, 0x53,
	0x7B, 0x38, 0x0D, 0x25, 0x22, 0x18, 0x0D, 0x07, 0x03, 0x06, 0x23, 0x06,
	0x35, 0x28, 0x29, 0x36, 0x0B, 0x0A, 0x3F, 0x53, 0x73, 0x3B, 0x18, 0x2A,
	0x3D, 0x11, 0x55, 0x50, 0x18, 0x07, 0x0E, 0x5C, 0x2F, 0x04, 0x2F, 0x10,
	0x01, 0x32, 0x5D, 0x0F, 0x69, 0x25, 0x37, 0x5E, 0x06, 0x0E, 0x0B, 0x27,
	0x0D, 0x08, 0x70, 0x5B, 0x0F, 0x41, 0x00, 0x2A, 0x1E, 0x13, 0x05, 0x12,
	0x15, 0x03, 0x07, 0x3A, 0x2E, 0x72, 0x21, 0x38, 0x5F, 0x58, 0x35, 0x20,
	0x37, 0x57, 0x3C, 0x11, 0x5F, 0x19, 0x09, 0x5B, 0x30, 0x1A, 0x0A, 0x1C,
	0x3A, 0x3B, 0x38, 0x39, 0x41, 0x26, 0x06, 0x21, 0x16, 0x2A, 0x09, 0x2B,
	0x2E, 0x08, 0x0F, 0x0D, 0x26, 0x23, 0x04, 0x36, 0x3C, 0x7B, 0x47, 0x2A,
	0x06, 0x25, 0x26, 0x0A, 0x1B, 0x24, 0x23, 0x35, 0x0F, 0x14, 0x5D, 0x18,
	0x07, 0x3A, 0x54, 0x02, 0x1D, 0x06, 0x1A, 0x17, 0x45, 0x44, 0x2B, 0x00,
	0x38, 0x17, 0x0E, 0x00, 0x16, 0x2D, 0x01, 0x5D, 0x35, 0x23, 0x0B, 0x45,
	0x1D, 0x33, 0x1F, 0x09, 0x1B, 0x00, 0x6D, 0x03, 0x26, 0x58, 0x39, 0x75,
	0x55, 0x37, 0x5F, 0x2C, 0x7B, 0x54, 0x29, 0x5B, 0x5C, 0x07, 0x5B, 0x4E,
	0x5F, 0x0F, 0x71, 0x03, 0x4E, 0x58, 0x1B, 0x05, 0x43, 0x54, 0x1D, 0x13,
	0x0C, 0x0E, 0x51, 0x17, 0x40, 0x3A, 0x5E, 0x2C, 0x1F, 0x13, 0x1B, 0x43,
	0x37, 0x14, 0x32, 0x23, 0x1E, 0x2B, 0x1D, 0x1C, 0x0F, 0x5B, 0x00, 0x5A,
	0x1B, 0x27, 0x14, 0x18, 0x5C, 0x1D, 0x3A, 0x5D, 0x11, 0x34, 0x0D, 0x16,
	0x27, 0x13, 0x25, 0x3F, 0x31, 0x2B, 0x00, 0x26, 0x3B, 0x05, 0x54, 0x06,
	0x07, 0x12, 0x7B, 0x58, 0x26, 0x29, 0x32, 0x28, 0x3E, 0x1B, 0x01, 0x1E,
	0x69, 0x2E, 0x14, 0x04, 0x29, 0x05, 0x00, 0x52, 0x04, 0x1D, 0x3A, 0x1B,
	0x0D, 0x17, 0x2F, 0x14, 0x05, 0x27, 0x0A, 0x3B, 0x01, 0x18, 0x2B, 0x45,
	0x1C, 0x1A, 0x3B, 0x18, 0x2F, 0x5A, 0x2A, 0x1B, 0x0D, 0x23, 0x2A, 0x26,
	0x2A, 0x0C, 0x3A, 0x01, 0x30, 0x5C, 0x24, 0x00, 0x02, 0x3A, 0x20, 0x32,
	0x17, 0x13, 0x71, 0x15, 0x0A, 0x5C, 0x26, 0x77, 0x16, 0x20, 0x5D, 0x5C,
	0x31, 0x5E, 0x0F, 0x56, 0x39, 0x37, 0x21, 0x2F, 0x16, 0x3D, 0x7A, 0x19,
	0x15, 0x2B, 0x19, 0x16, 0x03, 0x0C, 0x17, 0x38, 0x38, 0x15, 0x54, 0x00,
	0x0F, 0x70, 0x24, 0x4A, 0x01, 0x03, 0x24, 0x47, 0x55, 0x01, 0x2F, 0x08,
	0x0F, 0x39, 0x3B, 0x26, 0x76, 0x00, 0x4A, 0x5B, 0x2F, 0x0B, 0x19, 0x3B,
	0x3D, 0x40, 0x05, 0x1F, 0x0C, 0x59, 0x29, 0x20, 0x26, 0x23, 0x2A, 0x2A,
	0x69, 0x01, 0x11, 0x20, 0x52, 0x74, 0x3B, 0x39, 0x5B, 0x11, 0x2A, 0x55,
	0x18, 0x02, 0x3E, 0x1B, 0x04, 0x37, 0x1E, 0x5E, 0x05, 0x09, 0x31, 0x34,
	0x0C, 0x35, 0x3D, 0x27, 0x0B, 0x22, 0x7B, 0x2F, 0x50, 0x25, 0x44, 0x24,
	0x14, 0x17, 0x06, 0x18, 0x06, 0x3E, 0x30, 0x5F, 0x2C, 0x10, 0x21, 0x0E,
	0x25, 0x5B, 0x0D, 0x04, 0x27, 0x2C, 0x2C, 0x07, 0x09, 0x10, 0x05, 0x01,
	0x2B, 0x2B, 0x02, 0x06, 0x0F, 0x0D, 0x1D, 0x26, 0x3A, 0x27, 0x24, 0x55,
	0x27, 0x1C, 0x24, 0x2E, 0x0D, 0x15, 0x2D, 0x52, 0x24, 0x28, 0x0A, 0x2B,
	0x58, 0x1A, 0x43, 0x50, 0x2D, 0x3E, 0x0E, 0x34, 0x4A, 0x19, 0x5E, 0x00,
	0x00, 0x59, 0x39, 0x52, 0x28, 0x35, 0x23, 0x1C, 0x3A, 0x14, 0x39, 0x0A,
	0x36, 0x3B, 0x7B, 0x55, 0x36, 0x37, 0x26, 0x30, 0x58, 0x31, 0x21, 0x18,
	0x37, 0x26, 0x25, 0x0D, 0x1C, 0x75, 0x18, 0x29, 0x5A, 0x08, 0x13, 0x3E,
	0x12, 0x2B, 0x44, 0x7A, 0x28, 0x0A, 0x20, 0x1C, 0x17, 0x5C, 0x1B, 0x2A,
	0x1C, 0x01, 0x55, 0x08, 0x37, 0x3F, 0x05, 0x06, 0x27, 0x07, 0x1E, 0x2F,
	0x26, 0x38, 0x28, 0x04, 0x6D, 0x0A, 0x23, 0x2F, 0x32, 0x12, 0x1C, 0x36,
	0x0F, 0x38, 0x7B, 0x21, 0x19, 0x05, 0x5C, 0x34, 0x18, 0x3B, 0x23, 0x39,
	0x0A, 0x1D, 0x4E, 0x58, 0x20, 0x38, 0x35, 0x25, 0x2C, 0x23, 0x33, 0x58,
	0x04, 0x1F, 0x09, 0x72, 0x15, 0x07, 0x3C, 0x20, 0x2F, 0x59, 0x16, 0x58,
	0x13, 0x11, 0x29, 0x05, 0x16, 0x5B, 0x29, 0x2E, 0x36, 0x20, 0x1F, 0x37,
	0x58, 0x2E, 0x2C, 0x1D, 0x71, 0x2D, 0x53, 0x07, 0x1D, 0x06, 0x05, 0x37,
	0x25, 0x44, 0x77, 0x2F, 0x23, 0x59, 0x1D, 0x14, 0x1C, 0x34, 0x3F, 0x29,
	0x2B, 0x04, 0x3B, 0x1D, 0x18, 0x74, 0x24, 0x02, 0x5E, 0x06, 0x23, 0x38,
	0x09, 0x37, 0x2F, 0x25, 0x5A, 0x09, 0x17, 0x5B, 0x33, 0x1C, 0x58, 0x0A,
	0x1A, 0x29, 0x25, 0x23, 0x2B, 0x01, 0x13, 0x22, 0x05, 0x5D, 0x3D, 0x69,
	0x02, 0x2E, 0x07, 0x18, 0x35, 0x3D, 0x08, 0x21, 0x58, 0x0D, 0x2B, 0x2A,
	0x1F, 0x27, 0x07, 0x3E, 0x59, 0x5D, 0x23, 0x0B, 0x02, 0x0D, 0x5B, 0x07,
	0x11, 0x55, 0x4A, 0x20, 0x2E, 0x75, 0x25, 0x30, 0x06, 0x1A, 0x69, 0x27,
	0x37, 0x19, 0x20, 0x00, 0x55, 0x00, 0x5B, 0x2A, 0x1B, 0x2D, 0x14, 0x29,
	0x21, 0x69, 0x3E, 0x15, 0x0C, 0x33, 0x76, 0x00, 0x16, 0x3D, 0x1B, 0x14,
	0x3B, 0x0D, 0x5F, 0x0D, 0x21, 0x15, 0x30, 0x58, 0x27, 0x2B, 0x3B, 0x05,
	0x19, 0x3F, 0x13, 0x47, 0x25, 0x05, 0x3D, 0x0A, 0x5C, 0x3B, 0x02, 0x3E,
	0x75, 0x23, 0x23, 0x25, 0x2A, 0x3B, 0x08, 0x19, 0x41, 0x02, 0x28, 0x00,
	0x0F, 0x22, 0x25, 0x23, 0x3B, 0x11, 0x03, 0x5D, 0x13, 0x3C, 0x0A, 0x2D,
	0x59, 0x0B, 0x5C, 0x0F, 0x2F, 0x2F, 0x30, 0x09, 0x20, 0x01, 0x11, 0x34,
	0x18, 0x16, 0x07, 0x0C, 0x35, 0x59, 0x07, 0x56, 0x08, 0x35, 0x06, 0x2B,
	0x16, 0x25, 0x23, 0x0B, 0x34, 0x26, 0x1C, 0x6D, 0x2F, 0x2C, 0x39, 0x23,
	0x0A, 0x23, 0x0F, 0x59, 0x29, 0x07, 0x1C, 0x02, 0x04, 0x0F, 0x00, 0x5C,
	0x2E, 0x27, 0x52, 0x2C, 0x3A, 0x14, 0x21, 0x53, 0x35, 0x2B, 0x08, 0x3C,
	0x59, 0x69, 0x0F, 0x22, 0x59, 0x5B, 0x11, 0x2E, 0x14, 0x2F, 0x5A, 0x77,
	0x26, 0x51, 0x04, 0x2E, 0x6D, 0x3D, 0x36, 0x36, 0x23, 0x3B, 0x38, 0x08,
	0x3F, 0x1C, 0x1A, 0x24, 0x2A, 0x5A, 0x11, 0x7B, 0x35, 0x3B, 0x5B, 0x09,
	0x23, 0x26, 0x56, 0x0A, 0x3F, 0x76, 0x5B, 0x30, 0x1F, 0x33, 0x6D, 0x3F,
	0x28, 0x20, 0x39, 0x70, 0x2D, 0x0C, 0x1E, 0x02, 0x2A, 0x14, 0x55, 0x41,
	0x18, 0x72, 0x5E, 0x11, 0x0D, 0x0D, 0x1B, 0x1D, 0x36, 0x22, 0x03, 0x71,
	0x1B, 0x25, 0x3C, 0x06, 0x00, 0x19, 0x30, 0x0D, 0x00, 0x36, 0x47, 0x29,
	0x41, 0x29, 0x18, 0x16, 0x50, 0x0B, 0x13, 0x03, 0x18, 0x0B, 0x2F, 0x2A,
	0x0D, 0x05, 0x31, 0x0C, 0x2A, 0x77, 0x26, 0x2A, 0x36, 0x08, 0x70, 0x3E,
	0x3B, 0x56, 0x2F, 0x35, 0x38, 0x06, 0x0C, 0x07, 0x26, 0x43, 0x2C, 0x09,
	0x5C, 0x0D, 0x1E, 0x14, 0x23, 0x3B, 0x29, 0x08, 0x57, 0x23, 0x2E, 0x76,
	0x26, 0x27, 0x24, 0x40, 0x36, 0x14, 0x38, 0x0C, 0x00, 0x77, 0x0B, 0x20,
	0x18, 0x5C, 0x0D, 0x0B, 0x16, 0x38, 0x1B, 0x2A, 0x38, 0x2F, 0x27, 0x33,
	0x27, 0x5F, 0x02, 0x17, 0x0F, 0x06, 0x0F, 0x03, 0x1E, 0x29, 0x6D, 0x3C,
	0x17, 0x2A, 0x2D, 0x74, 0x1A, 0x4E, 0x41, 0x24, 0x0F, 0x54, 0x0D, 0x02,
	0x59, 0x2B, 0x3A, 0x2C, 0x2A, 0x44, 0x26, 0x5D, 0x3B, 0x1C, 0x5B, 0x74,
	0x2F, 0x39, 0x01, 0x3C, 0x35, 0x0B, 0x4A, 0x03, 0x3C, 0x30, 0x00, 0x59,
	0x0D, 0x0A, 0x2A, 0x0E, 0x35, 0x0C, 0x5D, 0x27, 0x5A, 0x37, 0x34, 0x3F,
	0x10, 0x15, 0x31, 0x18, 0x22, 0x2C, 0x03, 0x28, 0x58, 0x07, 0x26, 0x5A,
	0x39, 0x3E, 0x1D, 0x70, 0x28, 0x3B, 0x26, 0x53, 0x23, 0x5E, 0x51, 0x5D,
	0x5D, 0x23, 0x3B, 0x12, 0x00, 0x2F, 0x11, 0x2D, 0x59, 0x1C, 0x5F, 0x7B,
	0x04, 0x0D, 0x58, 0x1D, 0x76, 0x08, 0x51, 0x59, 0x02, 0x1B, 0x5F, 0x27,
	0x5A, 0x2F, 0x24, 0x58, 0x06, 0x37, 0x3B, 0x38, 0x23, 0x50, 0x04, 0x20,
	0x71, 0x05, 0x09, 0x02, 0x2F, 0x1A, 0x16, 0x13, 0x03, 0x1B, 0x76, 0x39,
	0x11, 0x59, 0x5E, 0x05, 0x3D, 0x05, 0x5C, 0x05, 0x32, 0x09, 0x0B, 0x0F,
	0x32, 0x04, 0x1C, 0x07, 0x04, 0x0C, 0x09, 0x28, 0x04, 0x41, 0x04, 0x0D,
	0x05, 0x05, 0x3F, 0x2C, 0x38, 0x58, 0x58, 0x07, 0x3B, 0x24, 0x59, 0x25,
	0x1F, 0x1A, 0x23, 0x5F, 0x39, 0x20, 0x3B, 0x24, 0x3B, 0x05, 0x5D, 0x5D,
	0x37, 0x5E, 0x05, 0x3B, 0x25, 0x6D, 0x01, 0x4E, 0x18, 0x29, 0x26, 0x55,
	0x51, 0x26, 0x26, 0x00, 0x0F, 0x53, 0x41, 0x01, 0x69, 0x06, 0x30, 0x59,
	0x29, 0x15, 0x18, 0x08, 0x5E, 0x3F, 0x23, 0x5D, 0x12, 0x21, 0x12, 0x2F,
	0x5F, 0x53, 0x29, 0x1F, 0x28, 0x54, 0x3B, 0x58, 0x28, 0x77, 0x21, 0x0E,
	0x24, 0x23, 0x36, 0x55, 0x4E, 0x02, 0x2A, 0x09, 0x15, 0x30, 0x58, 0x3D,
	0x25, 0x18, 0x55, 0x2A, 0x2C, 0x2A, 0x00, 0x36, 0x18, 0x3C, 0x29, 0x24,
	0x59, 0x02, 0x08, 0x6D, 0x54, 0x04, 0x14, 0x20, 0x0F, 0x24, 0x0A, 0x20,
	0x26, 0x73, 0x34, 0x2A, 0x0D, 0x0F, 0x0A, 0x27, 0x0C, 0x41, 0x29, 0x27,
	0x43, 0x33, 0x21, 0x06, 0x0E, 0x24, 0x59, 0x5A, 0x31, 0x20, 0x21, 0x2B,
	0x3D, 0x0D, 0x75, 0x54, 0x26, 0x59, 0x02, 0x25, 0x3A, 0x03, 0x1C, 0x0A,
	0x14, 0x43, 0x24, 0x02, 0x5C, 0x35, 0x5D, 0x27, 0x25, 0x32, 0x77, 0x3F,
	0x2C, 0x34, 0x3F, 0x21, 0x0F, 0x20, 0x20, 0x0F, 0x00, 0x43, 0x25, 0x58,
	0x02, 0x10, 0x1A, 0x3B, 0x0A, 0x32, 0x09, 0x2E, 0x39, 0x41, 0x0D, 0x31,
	0x3E, 0x05, 0x3F, 0x1D, 0x74, 0x47, 0x25, 0x41, 0x3A, 0x77, 0x0B, 0x2B,
	0x1B, 0x38, 0x1A, 0x2B, 0x50, 0x3A, 0x2F, 0x04, 0x5F, 0x19, 0x1E, 0x33,
	0x0F, 0x3D, 0x2F, 0x37, 0x2A, 0x2E, 0x16, 0x26, 0x28, 0x09, 0x2E, 0x23,
	0x35, 0x3E, 0x2C, 0x71, 0x28, 0x03, 0x3F, 0x3C, 0x14, 0x3E, 0x39, 0x5B,
	0x2C, 0x70, 0x27, 0x2D, 0x1F, 0x04, 0x36, 0x0F, 0x2E, 0x17, 0x44, 0x1B,
	0x47, 0x17, 0x1C, 0x5F, 0x28, 0x0E, 0x36, 0x08, 0x04, 0x14, 0x07, 0x2E,
	0x00, 0x1D, 0x15, 0x18, 0x16, 0x04, 0x53, 0x73, 0x39, 0x11, 0x57, 0x1C,
	0x33, 0x2A, 0x57, 0x5B, 0x0C, 0x17, 0x24, 0x50, 0x5B, 0x07, 0x05, 0x55,
	0x55, 0x56, 0x2C, 0x2E, 0x34, 0x51, 0x08, 0x2A, 0x73, 0x0A, 0x2F, 0x3C,
	0x2D, 0x69, 0x0E, 0x57, 0x56, 0x12, 0x07, 0x21, 0x03, 0x0A, 0x27, 0x72,
	0x2E, 0x20, 0x24, 0x02, 0x09, 0x15, 0x09, 0x3C, 0x33, 0x10, 0x1D, 0x58,
	0x37, 0x2D, 0x09, 0x22, 0x13, 0x3C, 0x08, 0x01, 0x2D, 0x07, 0x3B, 0x1F,
	0x69, 0x3C, 0x2C, 0x1A, 0x05, 0x38, 0x2D, 0x13, 0x2C, 0x3C, 0x0C, 0x16,
	0x2D, 0x45, 0x3F, 0x0A, 0x3A, 0x03, 0x5E, 0x32, 0x35, 0x5B, 0x17, 0x04,
	0x3E, 0x00, 0x16, 0x09, 0x16, 0x53, 0x14, 0x5F, 0x35, 0x1B, 0x3A, 0x0F,
	0x09, 0x29, 0x41, 0x5C, 0x01, 0x24, 0x3B, 0x41, 0x2C, 0x27, 0x54, 0x0F,
	0x28, 0x07, 0x2B, 0x2D, 0x11, 0x01, 0x0C, 0x38, 0x2D, 0x53, 0x34, 0x07,
	0x7B, 0x39, 0x24, 0x3A, 0x3E, 0x12, 0x15, 0x15, 0x08, 0x3F, 0x01, 0x08,
	0x2E, 0x21, 0x07, 0x0F, 0x55, 0x11, 0x5D, 0x2E, 0x31, 0x20, 0x05, 0x3F,
	0x02, 0x07, 0x43, 0x26, 0x1C, 0x3F, 0x72, 0x0E, 0x25, 0x2F, 0x0A, 0x36,
	0x07, 0x39, 0x26, 0x13, 0x2F, 0x5A, 0x57, 0x1A, 0x1B, 0x06, 0x23, 0x26,
	0x25, 0x19, 0x29, 0x35, 0x59, 0x5D, 0x59, 0x14, 0x36, 0x28, 0x0D, 0x1A,
	0x69, 0x0F, 0x3B, 0x26, 0x0D, 0x0A, 0x1B, 0x09, 0x3E, 0x13, 0x75, 0x07,
	0x18, 0x2A, 0x3F, 0x6D, 0x54, 0x0F, 0x5A, 0x27, 0x69, 0x0E, 0x0A, 0x03,
	0x26, 0x7B, 0x3F, 0x03, 0x39, 0x3A, 0x31, 0x00, 0x0A, 0x06, 0x40, 0x26,
	0x05, 0x31, 0x22, 0x05, 0x69, 0x26, 0x13, 0x02, 0x2A, 0x69, 0x2F, 0x17,
	0x25, 0x3A, 0x12, 0x19, 0x04, 0x20, 0x0D, 0x06, 0x03, 0x16, 0x16, 0x3E,
	0x26, 0x14, 0x00, 0x1C, 0x3F, 0x18, 0x28, 0x0F, 0x1E, 0x12, 0x77, 0x2E,
	0x2B, 0x3D, 0x52, 0x06, 0x34, 0x50, 0x5C, 0x2A, 0x2C, 0x59, 0x0D, 0x1A,
	0x13, 0x11, 0x18, 0x35, 0x1D, 0x5F, 0x34, 0x16, 0x34, 0x1A, 0x24, 0x17,
	0x39, 0x00, 0x1D, 0x25, 0x2E, 0x21, 0x59, 0x3F, 0x06, 0x03, 0x01, 0x28,
	0x27, 0x01, 0x2E, 0x3F, 0x09, 0x3B, 0x59, 0x33, 0x2A, 0x31, 0x5F, 0x0F,
	0x18, 0x1C, 0x15, 0x5E, 0x06, 0x13, 0x3D, 0x33, 0x41, 0x5B, 0x25, 0x01,
	0x07, 0x04, 0x12, 0x06, 0x3F, 0x34, 0x2C, 0x27, 0x2C, 0x1F, 0x2A, 0x5E,
	0x5E, 0x07, 0x06, 0x39, 0x56, 0x44, 0x31, 0x24, 0x22, 0x0F, 0x27, 0x04,
	0x39, 0x0D, 0x0D, 0x5F, 0x07, 0x5A, 0x02, 0x20, 0x44, 0x11, 0x19, 0x17,
	0x03, 0x0A, 0x7B, 0x1C, 0x13, 0x41, 0x0A, 0x27, 0x06, 0x55, 0x22, 0x33,
	0x21, 0x06, 0x2F, 0x24, 0x18, 0x7A, 0x22, 0x1B, 0x29, 0x58, 0x2B, 0x02,
	0x19, 0x5A, 0x1A, 0x1B, 0x27, 0x53, 0x2B, 0x07, 0x70, 0x07, 0x34, 0x56,
	0x1D, 0x34, 0x1B, 0x33, 0x24, 0x20, 0x35, 0x55, 0x0A, 0x2F, 0x39, 0x2B,
	0x38, 0x20, 0x5D, 0x0C, 0x20, 0x1B, 0x28, 0x07, 0x1F, 0x26, 0x3E, 0x28,
	0x28, 0x0E, 0x38, 0x14, 0x2C, 0x5A, 0x2D, 0x36, 0x38, 0x1B, 0x56, 0x25,
	0x1B, 0x1C, 0x0C, 0x5F, 0x1C, 0x2F, 0x36, 0x05, 0x08, 0x53, 0x21, 0x1F,
	0x09, 0x02, 0x3C, 0x01, 0x1C, 0x32, 0x1F, 0x44, 0x12, 0x59, 0x17, 0x16,
	0x53, 0x1A, 0x5B, 0x4A, 0x57, 0x0F, 0x0E, 0x43, 0x23, 0x39, 0x3A, 0x31,
	0x15, 0x1B, 0x3A, 0x22, 0x01, 0x2D, 0x16, 0x17, 0x5E, 0x13, 0x3F, 0x3B,
	0x3A, 0x03, 0x06, 0x3E, 0x1B, 0x06, 0x25, 0x29, 0x3F, 0x0E, 0x0D, 0x12,
	0x3B, 0x20, 0x19, 0x26, 0x0C, 0x36, 0x00, 0x17, 0x07, 0x3E, 0x33, 0x0E,
	0x36, 0x37, 0x1A, 0x0A, 0x29, 0x26, 0x3A, 0x5F, 0x29, 0x1D, 0x2A, 0x06,
	0x2F, 0x09, 0x02, 0x07, 0x1B, 0x38, 0x04, 0x2F, 0x0F, 0x1B, 0x5B, 0x0D,
	0x1C, 0x4A, 0x18, 0x33, 0x10, 0x43, 0x2A, 0x22, 0x1E, 0x05, 0x2B, 0x33,
	0x41, 0x24, 0x09, 0x39, 0x13, 0x5E, 0x0F, 0x69, 0x2D, 0x39, 0x2F, 0x0A,
	0x12, 0x20, 0x19, 0x00, 0x40, 0x1B, 0x14, 0x18, 0x3D, 0x05, 0x38, 0x05,
	0x51, 0x45, 0x38, 0x38, 0x20, 0x08, 0x34, 0x29, 0x24, 0x22, 0x0E, 0x23,
	0x1B, 0x06, 0x28, 0x03, 0x07, 0x27, 0x07, 0x3B, 0x2F, 0x3F, 0x3F, 0x16,
	0x27, 0x22, 0x2B, 0x20, 0x0D, 0x2E, 0x1B, 0x09, 0x5C, 0x08, 0x29, 0x12,
	0x3C, 0x0C, 0x2B, 0x5F, 0x39, 0x05, 0x40, 0x71, 0x47, 0x56, 0x25, 0x1E,
	0x13, 0x09, 0x24, 0x23, 0x22, 0x74, 0x2A, 0x16, 0x1F, 0x1D, 0x0A, 0x5B,
	0x34, 0x3E, 0x02, 0x2E, 0x3A, 0x56, 0x3B, 0x3C, 0x2D, 0x25, 0x54, 0x36,
	0x19, 0x74, 0x5F, 0x0B, 0x3D, 0x01, 0x16, 0x3A, 0x51, 0x3C, 0x01, 0x7B,
	0x0A, 0x39, 0x38, 0x32, 0x1A, 0x0B, 0x52, 0x1C, 0x21, 0x26, 0x1A, 0x2A,
	0x06, 0x28, 0x29, 0x29, 0x28, 0x1B, 0x0C, 0x0E, 0x22, 0x2F, 0x2C, 0x13,
	0x08, 0x55, 0x28, 0x2F, 0x3F, 0x11, 0x24, 0x2F, 0x29, 0x23, 0x73, 0x55,
	0x08, 0x36, 0x40, 0x2D, 0x2B, 0x13, 0x5B, 0x22, 0x0A, 0x1C, 0x39, 0x28,
	0x5D, 0x31, 0x5E, 0x22, 0x21, 0x3C, 0x17, 0x38, 0x35, 0x2A, 0x3E, 0x01,
	0x03, 0x04, 0x2A, 0x2E, 0x76, 0x05, 0x16, 0x18, 0x23, 0x35, 0x04, 0x0D,
	0x2B, 0x38, 0x26, 0x21, 0x56, 0x36, 0x08, 0x2B, 0x5C, 0x04, 0x2A, 0x39,
	0x01, 0x15, 0x36, 0x02, 0x53, 0x12, 0x18, 0x2B, 0x01, 0x3C, 0x25, 0x35,
	0x0C, 0x41, 0x2A, 0x04, 0x01, 0x28, 0x21, 0x53, 0x77, 0x27, 0x27, 0x37,
	0x01, 0x10, 0x38, 0x14, 0x07, 0x32, 0x70, 0x0F, 0x59, 0x27, 0x06, 0x26,
	0x25, 0x22, 0x1C, 0x2A, 0x2A, 0x24, 0x58, 0x45, 0x04, 0x38, 0x5B, 0x2F,
	0x58, 0x19, 0x2F, 0x23, 0x2C, 0x20, 0x5C, 0x06, 0x09, 0x09, 0x34, 0x28,
	0x12, 0x03, 0x00, 0x23, 0x5B, 0x2B, 0x24, 0x24, 0x5E, 0x25, 0x00, 0x35,
	0x2C, 0x24, 0x5E, 0x3B, 0x28, 0x28, 0x59, 0x5E, 0x26, 0x3E, 0x17, 0x09,
	0x5F, 0x29, 0x1F, 0x17, 0x08, 0x3F, 0x7A, 0x19, 0x07, 0x1F, 0x3F, 0x2A,
	0x35, 0x09, 0x25, 0x12, 0x34, 0x3E, 0x28, 0x5E, 0x05, 0x3A, 0x29, 0x14,
	0x03, 0x19, 0x33, 0x35, 0x03, 0x1F, 0x3D, 0x71, 0x5B, 0x03, 0x18, 0x29,
	0x06, 0x2E, 0x05, 0x3A, 0x5D, 0x27, 0x3E, 0x2D, 0x0F, 0x25, 0x73, 0x3F,
	0x2C, 0x39, 0x1D, 0x0F, 0x1C, 0x33, 0x41, 0x1A, 0x1B, 0x29, 0x35, 0x41,
	0x2E, 0x0C, 0x0D, 0x33, 0x08, 0x3F, 0x3B, 0x5C, 0x59, 0x18, 0x1D, 0x75,
	0x0D, 0x23, 0x5D, 0x26, 0x69, 0x1E, 0x06, 0x2B, 0x19, 0x14, 0x0F, 0x0D,
	0x3A, 0x58, 0x26, 0x1D, 0x07, 0x36, 0x12, 0x7A, 0x21, 0x56, 0x25, 0x3B,
	0x37, 0x3A, 0x0E, 0x08, 0x23, 0x3A, 0x1C, 0x19, 0x22, 0x09, 0x70, 0x3D,
	0x28, 0x3D, 0x19, 0x17, 0x38, 0x4A, 0x19, 0x26, 0x31, 0x54, 0x2F, 0x09,
	0x01, 0x73, 0x0B, 0x4E, 0x1F, 0x0D, 0x12, 0x3D, 0x34, 0x45, 0x04, 0x74,
	0x08, 0x09, 0x25, 0x05, 0x2F, 0x5F, 0x37, 0x19, 0x5B, 0x24, 0x22, 0x0E,
	0x18, 0x1C, 0x32, 0x1C, 0x39, 0x34, 0x59, 0x2B, 0x55, 0x24, 0x5F, 0x5F,
	0x00, 0x5E, 0x4E, 0x39, 0x24, 0x30, 0x0B, 0x39, 0x34, 0x0A, 0x70, 0x3F,
	0x57, 0x09, 0x5D, 0x36, 0x0B, 0x56, 0x58, 0x24, 0x3B, 0x2D, 0x57, 0x39,
	0x2F, 0x2F, 0x21, 0x05, 0x00, 0x2F, 0x35, 0x54, 0x52, 0x2A, 0x5E, 0x73,
	0x16, 0x07, 0x1F, 0x44, 0x0C, 0x1C, 0x2A, 0x0B, 0x09, 0x35, 0x16, 0x11,
	0x1E, 0x44, 0x20, 0x21, 0x51, 0x5E, 0x3F, 0x11, 0x2F, 0x3B, 0x56, 0x03,
	0x32, 0x5D, 0x57, 0x37, 0x2E, 0x09, 0x26, 0x0F, 0x2B, 0x3A, 0x72, 0x3D,
	0x51, 0x5A, 0x0D, 0x70, 0x3E, 0x2C, 0x56, 0x24, 0x18, 0x01, 0x16, 0x5B,
	0x18, 0x25, 0x5F, 0x36, 0x59, 0x01, 0x07, 0x08, 0x24, 0x3B, 0x1D, 0x18,
	0x47, 0x22, 0x1C, 0x40, 0x14, 0x43, 0x17, 0x3C, 0x3D, 0x0D, 0x0A, 0x04,
	0x09, 0x23, 0x6D, 0x34, 0x0E, 0x20, 0x00, 0x0D, 0x3A, 0x16, 0x1A, 0x08,
	0x09, 0x5B, 0x57, 0x0C, 0x3A, 0x01, 0x19, 0x24, 0x58, 0x08, 0x25, 0x29,
	0x11, 0x2A, 0x02, 0x1B, 0x5C, 0x10, 0x3B, 0x2F, 0x21, 0x09, 0x27, 0x01,
	0x31, 0x2D, 0x55, 0x13, 0x45, 0x2F, 0x15, 0x43, 0x26, 0x5A, 0x31, 0x08,
	0x08, 0x09, 0x25, 0x31, 0x77, 0x27, 0x18, 0x56, 0x25, 0x2A, 0x08, 0x56,
	0x1C, 0x08, 0x7A, 0x04, 0x19, 0x1C, 0x0D, 0x70, 0x27, 0x53, 0x34, 0x29,
	0x72, 0x5C, 0x0F, 0x36, 0x2F, 0x31, 0x2A, 0x22, 0x04, 0x31, 0x2A, 0x2F,
	0x0E, 0x36, 0x26, 0x70, 0x2F, 0x20, 0x21, 0x0A, 0x17, 0x1E, 0x2B, 0x2F,
	0x29, 0x1A, 0x28, 0x50, 0x0C, 0x1B, 0x7B, 0x3B, 0x58, 0x14, 0x5B, 0x10,
	0x22, 0x0C, 0x08, 0x3E, 0x70, 0x0A, 0x29, 0x3B, 0x59, 0x23, 0x55, 0x35,
	0x1D, 0x27, 0x0D, 0x06, 0x59, 0x2A, 0x19, 0x0C, 0x28, 0x50, 0x5F, 0x25,
	0x32, 0x16, 0x54, 0x57, 0x1C, 0x76, 0x0B, 0x00, 0x34, 0x1A, 0x76, 0x2B,
	0x2E, 0x1E, 0x02, 0x21, 0x2F, 0x06, 0x45, 0x33, 0x08, 0x05, 0x2B, 0x3C,
	0x58, 0x35, 0x04, 0x39, 0x5F, 0x24, 0x0C, 0x21, 0x57, 0x00, 0x2C, 0x31,
	0x5D, 0x14, 0x20, 0x39, 0x29, 0x58, 0x22, 0x06, 0x02, 0x18, 0x05, 0x58,
	0x0F, 0x32, 0x34, 0x23, 0x4A, 0x2C, 0x07, 0x2D, 0x2B, 0x31, 0x0D, 0x23,
	0x35, 0x09, 0x4A, 0x2C, 0x5D, 0x70, 0x07, 0x05, 0x5A, 0x0F, 0x73, 0x43,
	0x0E, 0x23, 0x3E, 0x27, 0x20, 0x35, 0x3C, 0x1B, 0x69, 0x14, 0x20, 0x45,
	0x58, 0x6D, 0x27, 0x0D, 0x45, 0x11, 0x29, 0x29, 0x51, 0x1A, 0x5C, 0x20,
	0x1F, 0x2E, 0x39, 0x53, 0x72, 0x03, 0x39, 0x56, 0x44, 0x24, 0x28, 0x08,
	0x09, 0x3D, 0x0B, 0x29, 0x53, 0x23, 0x0D, 0x35, 0x06, 0x2C, 0x26, 0x20,
	0x24, 0x59, 0x12, 0x21, 0x1A, 0x71, 0x09, 0x33, 0x5E, 0x59, 0x75, 0x3E,
	0x12, 0x03, 0x3C, 0x2A, 0x14, 0x08, 0x36, 0x08, 0x17, 0x2D, 0x0E, 0x2F,
	0x06, 0x28, 0x2D, 0x00, 0x1E, 0x38, 0x1A, 0x2E, 0x4E, 0x56, 0x5B, 0x17,
	0x29, 0x30, 0x2F, 0x59, 0x2F, 0x39, 0x30, 0x00, 0x1F, 0x70, 0x39, 0x24,
	0x57, 0x1A, 0x6D, 0x2B, 0x20, 0x38, 0x20, 0x12, 0x19, 0x18, 0x57, 0x08,
	0x77, 0x54, 0x0B, 0x28, 0x23, 0x09, 0x0D, 0x2E, 0x0A, 0x27, 0x14, 0x23,
	0x55, 0x20, 0x0E, 0x76, 0x16, 0x07, 0x3D, 0x38, 0x0A, 0x2D, 0x51, 0x2B,
	0x0D, 0x2D, 0x1F, 0x18, 0x19, 0x31, 0x04, 0x09, 0x2D, 0x3B, 0x1A, 0x2E,
	0x58, 0x17, 0x5B, 0x2C, 0x00, 0x5E, 0x08, 0x1E, 0x40, 0x72, 0x47, 0x09,
	0x00, 0x08, 0x0E, 0x16, 0x26, 0x2C, 0x38, 0x2B, 0x20, 0x31, 0x23, 0x24,
	0x06, 0x29, 0x04, 0x3E, 0x26, 0x31, 0x5B, 0x37, 0x07, 0x5D, 0x25, 0x34,
	0x35, 0x3C, 0x2A, 0x70, 0x5B, 0x4E, 0x58, 0x28, 0x6D, 0x3F, 0x05, 0x1B,
	0x0D, 0x2D, 0x1A, 0x58, 0x20, 0x13, 0x16, 0x27, 0x36, 0x28, 0x5B, 0x69,
	0x38, 0x13, 0x06, 0x5D, 0x13, 0x1C, 0x33, 0x1F, 0x39, 0x1A, 0x55, 0x0B,
	0x20, 0x2F, 0x35, 0x2D, 0x50, 0x3E, 0x2E, 0x0E, 0x47, 0x57, 0x1E, 0x2E,
	0x2B, 0x5F, 0x58, 0x34, 0x2A, 0x35, 0x24, 0x37, 0x00, 0x07, 0x29, 0x3C,
	0x18, 0x09, 0x1B, 0x37, 0x09, 0x10, 0x21, 0x24, 0x0D, 0x38, 0x59, 0x5F,
	0x2F, 0x13, 0x07, 0x38, 0x1E, 0x5A, 0x77, 0x59, 0x3B, 0x22, 0x05, 0x00,
	0x03, 0x2C, 0x5D, 0x5C, 0x11, 0x1C, 0x1B, 0x5D, 0x08, 0x28, 0x0E, 0x17,
	0x5B, 0x3F, 0x16, 0x1A, 0x0C, 0x24, 0x44, 0x27, 0x06, 0x11, 0x3A, 0x1C,
	0x17, 0x58, 0x1B, 0x59, 0x3C, 0x12, 0x26, 0x55, 0x1A, 0x20, 0x1B, 0x15,
	0x1B, 0x01, 0x1D, 0x15, 0x2B, 0x3B, 0x56, 0x25, 0x77, 0x38, 0x02, 0x03,
	0x29, 0x09, 0x1B, 0x38, 0x5D, 0x0C, 0x0F, 0x14, 0x52, 0x2D, 0x58, 0x73,
	0x20, 0x06, 0x3A, 0x5B, 0x70, 0x5C, 0x2B, 0x2D, 0x0C, 0x00, 0x5D, 0x25,
	0x36, 0x26, 0x7A, 0x2B, 0x26, 0x0B, 0x5D, 0x00, 0x2E, 0x24, 0x5E, 0x22,
	0x0B, 0x21, 0x17, 0x04, 0x1F, 0x00, 0x29, 0x58, 0x2D, 0x1C, 0x07, 0x05,
	0x08, 0x22, 0x3D, 0x11, 0x2B, 0x50, 0x38, 0x3A, 0x06, 0x3F, 0x14, 0x45,
	0x01, 0x1A, 0x1F, 0x14, 0x3D, 0x0A, 0x70, 0x27, 0x22, 0x07, 0x5F, 0x1B,
	0x04, 0x37, 0x39, 0x3F, 0x07, 0x3E, 0x2F, 0x5A, 0x0F, 0x6D, 0x59, 0x30,
	0x02, 0x1B, 0x31, 0x2A, 0x2D, 0x0F, 0x00, 0x76, 0x55, 0x1B, 0x2A, 0x5A,
	0x0F, 0x3C, 0x2E, 0x36, 0x08, 0x0D, 0x36, 0x09, 0x5A, 0x01, 0x26, 0x01,
	0x00, 0x02, 0x3A, 0x00, 0x07, 0x16, 0x57, 0x11, 0x16, 0x5D, 0x31, 0x41,
	0x3F, 0x23, 0x5E, 0x2E, 0x0B, 0x13, 0x6D, 0x2E, 0x36, 0x41, 0x5C, 0x2E,
	0x3A, 0x19, 0x02, 0x19, 0x16, 0x24, 0x55, 0x41, 0x00, 0x69, 0x24, 0x07,
	0x25, 0x5B, 0x1A, 0x1B, 0x16, 0x27, 0x04, 0x69, 0x09, 0x0E, 0x3C, 0x44,
	0x24, 0x5B, 0x22, 0x19, 0x00, 0x0D, 0x54, 0x13, 0x23, 0x21, 0x30, 0x58,
	0x24, 0x1C, 0x22, 0x7B, 0x00, 0x22, 0x1B, 0x0D, 0x03, 0x5B, 0x15, 0x29,
	0x11, 0x29, 0x26, 0x34, 0x3C, 0x28, 0x38, 0x24, 0x18, 0x03, 0x20, 0x74,
	0x54, 0x4A, 0x59, 0x2F, 0x0B, 0x16, 0x29, 0x57, 0x3F, 0x03, 0x18, 0x06,
	0x07, 0x5A, 0x2C, 0x55, 0x38, 0x56, 0x0D, 0x71, 0x03, 0x2E, 0x5E, 0x33,
	0x09, 0x3E, 0x13, 0x0F, 0x33, 0x28, 0x09, 0x0A, 0x28, 0x5C, 0x10, 0x22,
	0x18, 0x0C, 0x1C, 0x15, 0x0E, 0x03, 0x41, 0x27, 0x72, 0x22, 0x26, 0x5C,
	0x33, 0x74, 0x0D, 0x2E, 0x1A, 0x05, 0x26, 0x0F, 0x4E, 0x45, 0x3B, 0x10,
	0x3A, 0x09, 0x01, 0x3C, 0x13, 0x18, 0x17, 0x59, 0x03, 0x2C, 0x3A, 0x25,
	0x5C, 0x52, 0x7A, 0x23, 0x4A, 0x16, 0x2D, 0x2D, 0x3B, 0x1B, 0x2F, 0x18,
	0x0A, 0x2B, 0x51, 0x34, 0x11, 0x34, 0x25, 0x04, 0x29, 0x12, 0x01, 0x16,
	0x26, 0x23, 0x39, 0x20, 0x1F, 0x08, 0x07, 0x22, 0x15, 0x54, 0x2E, 0x3C,
	0x3D, 0x74, 0x03, 0x22, 0x3A, 0x3D, 0x25, 0x21, 0x33, 0x5F, 0x52, 0x10,
	0x3E, 0x58, 0x45, 0x12, 0x18, 0x0F, 0x02, 0x5E, 0x52, 0x09, 0x5F, 0x36,
	0x2B, 0x3D, 0x20, 0x24, 0x38, 0x3B, 0x0F, 0x33, 0x2B, 0x0C, 0x2D, 0x5B,
	0x7A, 0x19, 0x57, 0x17, 0x22, 0x12, 0x1E, 0x0C, 0x06, 0x09, 0x05, 0x18,
	0x2C, 0x05, 0x27, 0x24, 0x15, 0x59, 0x02, 0x00, 0x1B, 0x5D, 0x07, 0x2B,
	0x06, 0x11, 0x24, 0x1B, 0x57, 0x28, 0x27, 0x02, 0x06, 0x39, 0x1D, 0x0F,
	0x0D, 0x20, 0x56, 0x12, 0x32, 0x05, 0x22, 0x45, 0x2C, 0x0B, 0x35, 0x16,
	0x08, 0x2F, 0x07, 0x07, 0x58, 0x5A, 0x3A, 0x34, 0x1E, 0x55, 0x14, 0x44,
	0x12, 0x02, 0x19, 0x34, 0x26, 0x14, 0x5B, 0x0F, 0x38, 0x08, 0x34, 0x24,
	0x00, 0x59, 0x13, 0x33, 0x59, 0x2F, 0x2C, 0x1C, 0x1A, 0x1A, 0x39, 0x2D,
	0x05, 0x17, 0x24, 0x14, 0x29, 0x1F, 0x77, 0x22, 0x33, 0x03, 0x3D, 0x6D,
	0x3F, 0x53, 0x22, 0x0F, 0x24, 0x2A, 0x58, 0x2B, 0x40, 0x75, 0x5E, 0x26,
	0x22, 0x1B, 0x77, 0x03, 0x56, 0x21, 0x02, 0x75, 0x0E, 0x33, 0x28, 0x59,
	0x0B, 0x1E, 0x00, 0x3C, 0x32, 0x7B, 0x3A, 0x18, 0x19, 0x32, 0x18, 0x18,
	0x54, 0x57, 0x29, 0x27, 0x06, 0x0F, 0x22, 0x13, 0x0F, 0x3A, 0x06, 0x07,
	0x0F, 0x32, 0x5D, 0x08, 0x45, 0x0C, 0x69, 0x03, 0x04, 0x29, 0x04, 0x7A,
	0x34, 0x0C, 0x45, 0x2E, 0x01, 0x47, 0x2E, 0x1E, 0x3E, 0x06, 0x5F, 0x59,
	0x5B, 0x52, 0x30, 0x2B, 0x19, 0x1C, 0x5F, 0x38, 0x5C, 0x2C, 0x22, 0x04,
	0x30, 0x16, 0x34, 0x5F, 0x3B, 0x21, 0x15, 0x12, 0x2D, 0x32, 0x3B, 0x47,
	0x2F, 0x0A, 0x1C, 0x11, 0x55, 0x04, 0x0D, 0x5A, 0x17, 0x23, 0x59, 0x19,
	0x03, 0x26, 0x34, 0x03, 0x5D, 0x3F, 0x75, 0x15, 0x08, 0x36, 0x38, 0x36,
	0x0A, 0x30, 0x3D, 0x11, 0x3B, 0x35, 0x03, 0x1D, 0x22, 0x35, 0x01, 0x33,
	0x57, 0x1B, 0x07, 0x34, 0x56, 0x1A, 0x0F, 0x31, 0x25, 0x59, 0x26, 0x52,
	0x35, 0x1A, 0x4A, 0x28, 0x0D, 0x15, 0x3E, 0x10, 0x08, 0x52, 0x71, 0x23,
	0x2C, 0x2D, 0x12, 0x09, 0x5E, 0x34, 0x0B, 0x59, 0x2C, 0x01, 0x29, 0x57,
	0x04, 0x34, 0x5E, 0x22, 0x1D, 0x33, 0x04, 0x03, 0x16, 0x1D, 0x0D, 0x7B,
	0x0B, 0x06, 0x41, 0x23, 0x00, 0x1A, 0x02, 0x22, 0x3D, 0x0C, 0x03, 0x17,
	0x45, 0x2C, 0x03, 0x1F, 0x53, 0x17, 0x44, 0x76, 0x36, 0x22, 0x16, 0x23,
	0x16, 0x07, 0x2D, 0x41, 0x25, 0x6D, 0x1F, 0x27, 0x08, 0x05, 0x70, 0x43,
	0x16, 0x27, 0x44, 0x0E, 0x55, 0x07, 0x18, 0x52, 0x29, 0x27, 0x23, 0x0C,
	0x19, 0x27, 0x00, 0x4A, 0x1B, 0x58, 0x3A, 0x3C, 0x16, 0x21, 0x1B, 0x33,
	0x05, 0x50, 0x02, 0x40, 0x12, 0x47, 0x55, 0x37, 0x58, 0x06, 0x27, 0x36,
	0x59, 0x39, 0x28, 0x29, 0x51, 0x5A, 0x5C, 0x00, 0x1E, 0x04, 0x19, 0x1E,
	0x24, 0x1F, 0x2D, 0x37, 0x23, 0x75, 0x08, 0x0B, 0x5E, 0x25, 0x7A, 0x01,
	0x37, 0x0C, 0x1F, 0x0D, 0x18, 0x29, 0x2C, 0x3D, 0x14, 0x18, 0x0E, 0x14,
	0x1C, 0x0C, 0x15, 0x03, 0x2A, 0x06, 0x24, 0x3A, 0x37, 0x26, 0x5D, 0x28,
	0x2D, 0x59, 0x26, 0x5B, 0x0B, 0x25, 0x25, 0x1E, 0x23, 0x25, 0x2E, 0x35,
	0x21, 0x5F, 0x08, 0x1C, 0x54, 0x57, 0x3F, 0x2B, 0x19, 0x31, 0x58, 0x12,
	0x35, 0x25, 0x29, 0x0F, 0x20, 0x3A, 0x43, 0x24, 0x1F, 0x33, 0x14, 0x3B,
	0x53, 0x58, 0x02, 0x21, 0x24, 0x02, 0x1C, 0x31, 0x36, 0x34, 0x2B, 0x5C,
	0x20, 0x05, 0x09, 0x0B, 0x0D, 0x07, 0x04, 0x35, 0x56, 0x03, 0x53, 0x6D,
	0x34, 0x22, 0x5A, 0x0A, 0x3B, 0x5B, 0x52, 0x17, 0x1C, 0x69, 0x3B, 0x2C,
	0x02, 0x1F, 0x23, 0x34, 0x0F, 0x18, 0x02, 0x00, 0x21, 0x08, 0x37, 0x04,
	0x21, 0x5F, 0x04, 0x18, 0x31, 0x14, 0x15, 0x4A, 0x29, 0x28, 0x3A, 0x01,
	0x00, 0x36, 0x05, 0x32, 0x23, 0x15, 0x16, 0x2F, 0x21, 0x23, 0x20, 0x0B,
	0x1C, 0x28, 0x5C, 0x16, 0x3F, 0x07, 0x04, 0x24, 0x09, 0x21, 0x19, 0x2B,
	0x19, 0x26, 0x06, 0x26, 0x0D, 0x2B, 0x36, 0x23, 0x31, 0x30, 0x0E, 0x17,
	0x0B, 0x5D, 0x0F, 0x21, 0x28, 0x38, 0x12, 0x76, 0x03, 0x18, 0x41, 0x2F,
	0x2A, 0x35, 0x28, 0x05, 0x58, 0x07, 0x5F, 0x38, 0x5D, 0x1C, 0x06, 0x35,
	0x29, 0x22, 0x32, 0x6D, 0x5E, 0x10, 0x1A, 0x0F, 0x36, 0x3E, 0x56, 0x19,
	0x3F, 0x34, 0x5E, 0x16, 0x27, 0x09, 0x2B, 0x1A, 0x53, 0x38, 0x1E, 0x77,
	0x38, 0x56, 0x26, 0x08, 0x21, 0x2E, 0x23, 0x16, 0x28, 0x0E, 0x21, 0x0C,
	0x56, 0x32, 0x00, 0x36, 0x0B, 0x37, 0x03, 0x18, 0x1F, 0x59, 0x34, 0x5B,
	0x70, 0x58, 0x0C, 0x0F, 0x24, 0x1B, 0x36, 0x09, 0x5F, 0x19, 0x73, 0x06,
	0x15, 0x24, 0x5B, 0x2D, 0x27, 0x4E, 0x57, 0x53, 0x17, 0x1C, 0x59, 0x08,
	0x0C, 0x73, 0x00, 0x36, 0x3F, 0x28, 0x72, 0x06, 0x30, 0x58, 0x58, 0x11,
	0x0B, 0x08, 0x1E, 0x21, 0x1B, 0x3A, 0x15, 0x3C, 0x28, 0x37, 0x54, 0x04,
	0x21, 0x29, 0x00, 0x0D, 0x34, 0x56, 0x24, 0x70, 0x03, 0x17, 0x27, 0x3A,
	0x31, 0x0A, 0x03, 0x0A, 0x2A, 0x33, 0x04, 0x0A, 0x5B, 0x3A, 0x37, 0x38,
	0x09, 0x07, 0x29, 0x2B, 0x5B, 0x03, 0x45, 0x2D, 0x0B, 0x3A, 0x03, 0x57,
	0x27, 0x16, 0x54, 0x22, 0x1D, 0x0A, 0x3B, 0x2D, 0x36, 0x3B, 0x05, 0x2A,
	0x09, 0x50, 0x28, 0x33, 0x23, 0x34, 0x57, 0x1C, 0x5B, 0x12, 0x1E, 0x2F,
	0x0A, 0x52, 0x69, 0x20, 0x12, 0x06, 0x32, 0x2C, 0x14, 0x04, 0x28, 0x06,
	0x14, 0x2F, 0x2C, 0x18, 0x3E, 0x75, 0x35, 0x11, 0x34, 0x12, 0x72, 0x39,
	0x08, 0x16, 0x1D, 0x11, 0x0A, 0x30, 0x3E, 0x22, 0x15, 0x04, 0x18, 0x36,
	0x03, 0x0E, 0x18, 0x33, 0x3B, 0x24, 0x38, 0x3C, 0x31, 0x5F, 0x0C, 0x31,
	0x2B, 0x0E, 0x1B, 0x52, 0x6D, 0x25, 0x31, 0x28, 0x01, 0x08, 0x0E, 0x26,
	0x02, 0x13, 0x75, 0x5B, 0x4E, 0x07, 0x22, 0x2F, 0x27, 0x25, 0x25, 0x1B,
	0x36, 0x15, 0x2A, 0x2F, 0x3E, 0x14, 0x06, 0x2A, 0x01, 0x19, 0x35, 0x5C,
	0x37, 0x26, 0x0C, 0x16, 0x2E, 0x58, 0x0D, 0x05, 0x21, 0x00, 0x02, 0x25,
	0x03, 0x2F, 0x35, 0x34, 0x00, 0x24, 0x1A, 0x3B, 0x22, 0x1F, 0x26, 0x10,
	0x08, 0x25, 0x06, 0x0C, 0x34, 0x06, 0x58, 0x1E, 0x28, 0x25, 0x3D, 0x34,
	0x5B, 0x3E, 0x25, 0x03, 0x07, 0x14, 0x19, 0x0C, 0x18, 0x0B, 0x5F, 0x0E,
	0x77, 0x15, 0x2E, 0x3E, 0x1B, 0x0A, 0x0A, 0x0B, 0x27, 0x44, 0x12, 0x38,
	0x53, 0x39, 0x1C, 0x6D, 0x01, 0x07, 0x59, 0x44, 0x04, 0x2E, 0x4E, 0x2C,
	0x05, 0x27, 0x23, 0x04, 0x45, 0x26, 0x28, 0x26, 0x15, 0x26, 0x2A, 0x69,
	0x0F, 0x11, 0x1C, 0x0F, 0x3A, 0x36, 0x58, 0x22, 0x40, 0x6D, 0x54, 0x31,
	0x26, 0x52, 0x2C, 0x20, 0x0D, 0x41, 0x1C, 0x2D, 0x3C, 0x13, 0x25, 0x58,
	0x7A, 0x3C, 0x58, 0x04, 0x3B, 0x36, 0x25, 0x31, 0x5F, 0x24, 0x0F, 0x0B,
	0x29, 0x56, 0x2C, 0x28, 0x2D, 0x53, 0x16, 0x25, 0x33, 0x3B, 0x13, 0x26,
	0x1F, 0x1B, 0x1B, 0x17, 0x39, 0x3A, 0x12, 0x58, 0x0E, 0x25, 0x5E, 0x11,
	0x3B, 0x2D, 0x5B, 0x26, 0x14, 0x15, 0x0C, 0x00, 0x06, 0x31, 0x58, 0x26,
	0x45, 0x3A, 0x33, 0x59, 0x28, 0x0F, 0x00, 0x20, 0x2A, 0x27, 0x14, 0x3A,
	0x18, 0x54, 0x04, 0x07, 0x12, 0x26, 0x24, 0x1B, 0x0F, 0x03, 0x12, 0x01,
	0x25, 0x1B, 0x1C, 0x3A, 0x01, 0x4A, 0x34, 0x18, 0x06, 0x59, 0x38, 0x1C,
	0x01, 0x0F, 0x05, 0x0C, 0x29, 0x0F, 0x01, 0x16, 0x00, 0x0C, 0x09, 0x32,
	0x5E, 0x35, 0x3F, 0x25, 0x24, 0x16, 0x04, 0x2B, 0x18, 0x2F, 0x01, 0x36,
	0x2C, 0x5C, 0x0C, 0x1C, 0x19, 0x01, 0x5A, 0x17, 0x16, 0x06, 0x25, 0x08,
	0x73, 0x0F, 0x17, 0x5F, 0x0A, 0x09, 0x3D, 0x2F, 0x3A, 0x1C, 0x12, 0x0D,
	0x15, 0x27, 0x32, 0x73, 0x1A, 0x0E, 0x1A, 0x58, 0x0D, 0x5C, 0x0A, 0x01,
	0x19, 0x69, 0x0E, 0x05, 0x05, 0x59, 0x01, 0x22, 0x37, 0x5A, 0x0E, 0x24,
	0x05, 0x08, 0x14, 0x5D, 0x1A, 0x29, 0x13, 0x3A, 0x04, 0x15, 0x2E, 0x26,
	0x5E, 0x23, 0x1A, 0x36, 0x34, 0x24, 0x2D, 0x33, 0x1E, 0x02, 0x0B, 0x2E,
	0x36, 0x1C, 0x0C, 0x5F, 0x5D, 0x2D, 0x0B, 0x35, 0x09, 0x08, 0x00, 0x02,
	0x16, 0x36, 0x08, 0x20, 0x38, 0x12, 0x25, 0x5C, 0x73, 0x5C, 0x56, 0x1F,
	0x1C, 0x38, 0x03, 0x24, 0x20, 0x31, 0x37, 0x5C, 0x0C, 0x1D, 0x53, 0x21,
	0x0B, 0x50, 0x0A, 0x07, 0x7A, 0x29, 0x07, 0x17, 0x3D, 0x75, 0x2D, 0x12,
	0x02, 0x24, 0x16, 0x04, 0x36, 0x25, 0x11, 0x08, 0x1E, 0x57, 0x5A, 0x3F,
	0x24, 0x2A, 0x27, 0x1C, 0x3B, 0x74, 0x28, 0x22, 0x1B, 0x0D, 0x0B, 0x55,
	0x26, 0x37, 0x20, 0x15, 0x15, 0x23, 0x22, 0x44, 0x31, 0x43, 0x2D, 0x3A,
	0x0A, 0x2D, 0x03, 0x52, 0x1E, 0x20, 0x76, 0x06, 0x03, 0x09, 0x12, 0x01,
	0x36, 0x57, 0x21, 0x39, 0x26, 0x1B, 0x14, 0x24, 0x5D, 0x03, 0x2B, 0x26,
	0x3A, 0x06, 0x08, 0x16, 0x08, 0x57, 0x19, 0x74, 0x15, 0x35, 0x23, 0x11,
	0x20, 0x2A, 0x28, 0x1E, 0x5C, 0x2A, 0x36, 0x17, 0x3D, 0x28, 0x72, 0x26,
	0x27, 0x01, 0x18, 0x04, 0x3E, 0x0B, 0x45, 0x04, 0x36, 0x5E, 0x2B, 0x17,
	0x18, 0x04, 0x0B, 0x02, 0x59, 0x12, 0x75, 0x18, 0x15, 0x0A, 0x01, 0x23,
	0x35, 0x2D, 0x2B, 0x2E, 0x71, 0x1A, 0x50, 0x1F, 0x19, 0x7A, 0x3B, 0x59,
	0x19, 0x3C, 0x08, 0x26, 0x17, 0x26, 0x1F, 0x00, 0x1E, 0x59, 0x38, 0x40,
	0x04, 0x3F, 0x18, 0x39, 0x1C, 0x30, 0x1A, 0x29, 0x57, 0x5A, 0x32, 0x21,
	0x22, 0x06, 0x32, 0x20, 0x2E, 0x09, 0x3F, 0x58, 0x31, 0x20, 0x05, 0x07,
	0x13, 0x21, 0x2A, 0x08, 0x34, 0x1F, 0x74, 0x55, 0x14, 0x57, 0x0F, 0x2B,
	0x0D, 0x55, 0x22, 0x2D, 0x17, 0x02, 0x0F, 0x5D, 0x59, 0x75, 0x5C, 0x36,
	0x0B, 0x12, 0x14, 0x35, 0x2D, 0x27, 0x5A, 0x71, 0x3C, 0x58, 0x20, 0x19,
	0x0F, 0x39, 0x4A, 0x19, 0x59, 0x09, 0x5E, 0x59, 0x45, 0x5D, 0x77, 0x09,
	0x09, 0x45, 0x2A, 0x0D, 0x2A, 0x12, 0x1D, 0x2A, 0x7B, 0x0E, 0x39, 0x36,
	0x32, 0x33, 0x59, 0x06, 0x1D, 0x3A, 0x2F, 0x54, 0x4A, 0x5E, 0x1A, 0x34,
	0x06, 0x03, 0x5A, 0x08, 0x0E, 0x26, 0x03, 0x28, 0x1E, 0x6D, 0x43, 0x3B,
	0x0D, 0x11, 0x07, 0x3D, 0x09, 0x3D, 0x0F, 0x00, 0x5C, 0x05, 0x3B, 0x04,
	0x01, 0x5B, 0x0E, 0x18, 0x3A, 0x10, 0x00, 0x3B, 0x17, 0x21, 0x28, 0x39,
	0x37, 0x56, 0x5D, 0x26, 0x27, 0x50, 0x36, 0x13, 0x0F, 0x5C, 0x0E, 0x14,
	0x2A, 0x7A, 0x39, 0x2C, 0x01, 0x09, 0x23, 0x05, 0x58, 0x3E, 0x53, 0x18,
	0x35, 0x0F, 0x38, 0x5D, 0x27, 0x5F, 0x10, 0x00, 0x5F, 0x0C, 0x15, 0x0D,
	0x00, 0x23, 0x35, 0x3E, 0x2F, 0x59, 0x05, 0x7A, 0x0B, 0x14, 0x17, 0x0E,
	0x2A, 0x2D, 0x37, 0x0D, 0x5C, 0x20, 0x2B, 0x59, 0x2D, 0x53, 0x7B, 0x00,
	0x39, 0x2D, 0x00, 0x38, 0x54, 0x11, 0x5B, 0x44, 0x08, 0x0D, 0x22, 0x1A,
	0x21, 0x32, 0x43, 0x0F, 0x20, 0x12, 0x18, 0x35, 0x08, 0x16, 0x24, 0x34,
	0x00, 0x24, 0x36, 0x13, 0x2C, 0x1A, 0x59, 0x34, 0x02, 0x0D, 0x1E, 0x25,
	0x36, 0x05, 0x1A, 0x1F, 0x53, 0x0B, 0x5F, 0x72, 0x03, 0x12, 0x34, 0x5A,
	0x0F, 0x1E, 0x1B, 0x26, 0x05, 0x14, 0x1F, 0x0A, 0x1F, 0x00, 0x35, 0x15,
	0x20, 0x3F, 0x23, 0x33, 0x1A, 0x50, 0x09, 0x23, 0x33, 0x20, 0x4E, 0x01,
	0x26, 0x0C, 0x26, 0x52, 0x0D, 0x13, 0x2A, 0x55, 0x56, 0x57, 0x09, 0x32,
	0x47, 0x56, 0x00, 0x3D, 0x76, 0x08, 0x0D, 0x17, 0x13, 0x6D, 0x3B, 0x38,
	0x22, 0x09, 0x26, 0x0F, 0x2C, 0x36, 0x40, 0x31, 0x5C, 0x4E, 0x08, 0x39,
	0x0A, 0x27, 0x0C, 0x2C, 0x5B, 0x1A, 0x0F, 0x54, 0x17, 0x5E, 0x18, 0x1E,
	0x06, 0x02, 0x0D, 0x33, 0x5A, 0x14, 0x3E, 0x03, 0x2E, 0x22, 0x06, 0x3E,
	0x1A, 0x20, 0x3E, 0x4E, 0x20, 0x5E, 0x2D, 0x1A, 0x35, 0x28, 0x2E, 0x24,
	0x2D, 0x18, 0x5C, 0x1E, 0x2F, 0x23, 0x50, 0x3F, 0x3D, 0x15, 0x3E, 0x1B,
	0x2C, 0x05, 0x1A, 0x1E, 0x36, 0x37, 0x5A, 0x1B, 0x59, 0x04, 0x3D, 0x1A,
	0x7A, 0x1B, 0x23, 0x00, 0x12, 0x38, 0x5B, 0x04, 0x08, 0x0A, 0x3B, 0x43,
	0x33, 0x1C, 0x26, 0x71, 0x03, 0x39, 0x2F, 0x0D, 0x25, 0x15, 0x0A, 0x0F,
	0x2C, 0x0C, 0x1A, 0x35, 0x1B, 0x31, 0x71, 0x02, 0x59, 0x45, 0x53, 0x35,
	0x0B, 0x58, 0x0C, 0x00, 0x18, 0x5D, 0x36, 0x09, 0x11, 0x70, 0x5E, 0x55,
	0x07, 0x5F, 0x35, 0x36, 0x22, 0x38, 0x05, 0x70, 0x1D, 0x04, 0x3C, 0x21,
	0x33, 0x5F, 0x20, 0x59, 0x0E, 0x16, 0x5A, 0x28, 0x56, 0x07, 0x08, 0x5B,
	0x0B, 0x18, 0x38, 0x73, 0x16, 0x07, 0x1D, 0x00, 0x01, 0x1A, 0x35, 0x02,
	0x21, 0x01, 0x0A, 0x0D, 0x01, 0x20, 0x6D, 0x2F, 0x28, 0x38, 0x2D, 0x11,
	0x5E, 0x07, 0x5B, 0x12, 0x7A, 0x00, 0x58, 0x09, 0x38, 0x0D, 0x01, 0x37,
	0x2F, 0x07, 0x27, 0x3B, 0x55, 0x19, 0x06, 0x31, 0x23, 0x0E, 0x03, 0x5C,
	0x29, 0x0B, 0x15, 0x1D, 0x5B, 0x29, 0x01, 0x34, 0x17, 0x2C, 0x0F, 0x2E,
	0x39, 0x20, 0x1E, 0x06, 0x03, 0x1B, 0x03, 0x28, 0x07, 0x28, 0x19, 0x0F,
	0x1B, 0x6D, 0x21, 0x37, 0x2F, 0x2C, 0x74, 0x0E, 0x1B, 0x02, 0x08, 0x69,
	0x0B, 0x53, 0x29, 0x19, 0x34, 0x16, 0x12, 0x0B, 0x5F, 0x33, 0x38, 0x14,
	0x00, 0x40, 0x33, 0x1A, 0x31, 0x05, 0x3A, 0x1B, 0x19, 0x2E, 0x1F, 0x1D,
	0x1B, 0x3B, 0x00, 0x08, 0x03, 0x7B, 0x5E, 0x0B, 0x05, 0x5A, 0x08, 0x38,
	0x0D, 0x0B, 0x5E, 0x29, 0x1B, 0x0B, 0x04, 0x5F, 0x1B, 0x54, 0x08, 0x1F,
	0x44, 0x2C, 0x3D, 0x34, 0x1B, 0x3B, 0x37, 0x5E, 0x38, 0x2F, 0x53, 0x23,
	0x03, 0x35, 0x57, 0x1A, 0x7A, 0x47, 0x27, 0x19, 0x2E, 0x0A, 0x47, 0x27,
	0x16, 0x0E, 0x33, 0x23, 0x24, 0x3D, 0x24, 0x31, 0x3A, 0x0C, 0x0A, 0x53,
	0x04, 0x47, 0x56, 0x38, 0x18, 0x1B, 0x3A, 0x15, 0x2F, 0x08, 0x23, 0x3C,
	0x03, 0x03, 0x09, 0x20, 0x27, 0x03, 0x01, 0x53, 0x69, 0x25, 0x02, 0x36,
	0x32, 0x23, 0x0D, 0x04, 0x3E, 0x32, 0x2B, 0x55, 0x35, 0x0D, 0x02, 0x10,
	0x1E, 0x03, 0x29, 0x02, 0x33, 0x5A, 0x27, 0x28, 0x07, 0x00, 0x27, 0x0D,
	0x19, 0x5F, 0x0E, 0x34, 0x0A, 0x3F, 0x29, 0x1A, 0x06, 0x12, 0x3F, 0x3C,
	0x2A, 0x5D, 0x35, 0x1A, 0x38, 0x12, 0x08, 0x1B, 0x1B, 0x5F, 0x16, 0x5C,
	0x2A, 0x1A, 0x08, 0x32, 0x2D, 0x27, 0x0D, 0x1B, 0x76, 0x19, 0x35, 0x22,
	0x13, 0x27, 0x04, 0x37, 0x0A, 0x5D, 0x2D, 0x00, 0x51, 0x17, 0x0D, 0x77,
	0x34, 0x03, 0x5B, 0x32, 0x2A, 0x16, 0x04, 0x1E, 0x33, 0x76, 0x5A, 0x34,
	0x28, 0x2C, 0x37, 0x1C, 0x36, 0x41, 0x1A, 0x0C, 0x47, 0x08, 0x17, 0x06,
	0x28, 0x34, 0x2E, 0x0B, 0x5D, 0x15, 0x02, 0x0D, 0x3D, 0x2D, 0x30, 0x5D,
	0x38, 0x41, 0x22, 0x35, 0x3A, 0x52, 0x16, 0x00, 0x74, 0x2F, 0x51, 0x3E,
	0x53, 0x7A, 0x0A, 0x16, 0x3D, 0x19, 0x71, 0x00, 0x51, 0x22, 0x3E, 0x1B,
	0x54, 0x31, 0x37, 0x21, 0x35, 0x03, 0x23, 0x00, 0x1D, 0x37, 0x58, 0x23,
	0x2F, 0x40, 0x77, 0x5A, 0x10, 0x3C, 0x08, 0x0F, 0x19, 0x26, 0x0C, 0x40,
	0x12, 0x47, 0x11, 0x5F, 0x44, 0x37, 0x54, 0x4A, 0x07, 0x05, 0x75, 0x02,
	0x16, 0x41, 0x1F, 0x6D, 0x1E, 0x07, 0x05, 0x40, 0x15, 0x5B, 0x02, 0x14,
	0x31, 0x76, 0x3A, 0x0B, 0x25, 0x5F, 0x72, 0x07, 0x03, 0x3D, 0x53, 0x13,
	0x1C, 0x26, 0x21, 0x04, 0x08, 0x1E, 0x2D, 0x5F, 0x07, 0x0D, 0x1D, 0x58,
	0x25, 0x2E, 0x33, 0x24, 0x36, 0x22, 0x59, 0x24, 0x43, 0x34, 0x03, 0x19,
	0x36, 0x5C, 0x2A, 0x1C, 0x2D, 0x7A, 0x1D, 0x13, 0x0C, 0x5E, 0x71, 0x2D,
	0x22, 0x39, 0x1B, 0x07, 0x38, 0x39, 0x1C, 0x18, 0x38, 0x15, 0x2F, 0x1A,
	0x11, 0x20, 0x1D, 0x11, 0x36, 0x01, 0x27, 0x16, 0x04, 0x26, 0x5F, 0x06,
	0x29, 0x13, 0x1D, 0x12, 0x26, 0x16, 0x03, 0x23, 0x19, 0x74, 0x38, 0x10,
	0x03, 0x27, 0x15, 0x0E, 0x05, 0x14, 0x0D, 0x33, 0x15, 0x57, 0x3F, 0x28,
	0x14, 0x27, 0x2F, 0x39, 0x05, 0x03, 0x5D, 0x36, 0x0B, 0x2C, 0x16, 0x26,
	0x25, 0x5F, 0x3A, 0x76, 0x29, 0x2C, 0x01, 0x1A, 0x0F, 0x3A, 0x09, 0x06,
	0x27, 0x04, 0x14, 0x11, 0x2A, 0x19, 0x0B, 0x0E, 0x08, 0x08, 0x0F, 0x17,
	0x03, 0x13, 0x2C, 0x1C, 0x0F, 0x25, 0x57, 0x3B, 0x33, 0x18, 0x25, 0x03,
	0x41, 0x33, 0x05, 0x5A, 0x17, 0x57, 0x19, 0x2D, 0x07, 0x05, 0x5C, 0x5B,
	0x2A, 0x2A, 0x33, 0x5C, 0x0D, 0x05, 0x1A, 0x55, 0x1C, 0x38, 0x0D, 0x36,
	0x0D, 0x1F, 0x2F, 0x0E, 0x01, 0x1B, 0x57, 0x0E, 0x24, 0x07, 0x33, 0x1A,
	0x04, 0x17, 0x55, 0x28, 0x39, 0x1C, 0x25, 0x59, 0x13, 0x07, 0x3C, 0x16,
	0x18, 0x2B, 0x1F, 0x40, 0x0E, 0x5D, 0x2B, 0x0C, 0x40, 0x0F, 0x23, 0x28,
	0x0D, 0x26, 0x27, 0x5D, 0x25, 0x57, 0x07, 0x26, 0x43, 0x27, 0x57, 0x23,
	0x6D, 0x29, 0x09, 0x1A, 0x32, 0x17, 0x05, 0x55, 0x1A, 0x1F, 0x00, 0x1F,
	0x57, 0x20, 0x5A, 0x38, 0x28, 0x34, 0x3C, 0x1A, 0x6D, 0x07, 0x04, 0x5A,
	0x19, 0x2D, 0x2A, 0x38, 0x3E, 0x00, 0x16, 0x16, 0x39, 0x08, 0x1D, 0x7B,
	0x28, 0x19, 0x34, 0x2F, 0x77, 0x5B, 0x36, 0x38, 0x58, 0x73, 0x43, 0x24,
	0x2D, 0x2E, 0x17, 0x09, 0x50, 0x27, 0x18, 0x76, 0x19, 0x25, 0x37, 0x04,
	0x7A, 0x34, 0x12, 0x3F, 0x53, 0x2D, 0x09, 0x4A, 0x2B, 0x24, 0x73, 0x3F,
	0x1B, 0x0D, 0x33, 0x7B, 0x01, 0x31, 0x20, 0x0A, 0x14, 0x01, 0x59, 0x28,
	0x5B, 0x0A, 0x01, 0x15, 0x26, 0x53, 0x2B, 0x20, 0x30, 0x14, 0x3F, 0x24,
	0x22, 0x30, 0x08, 0x33, 0x03, 0x1F, 0x2C, 0x1F, 0x0A, 0x31, 0x3B, 0x52,
	0x04, 0x0E, 0x18, 0x05, 0x52, 0x29, 0x04, 0x07, 0x24, 0x00, 0x2B, 0x3B,
	0x74, 0x2D, 0x06, 0x2C, 0x58, 0x2C, 0x5F, 0x0A, 0x2B, 0x00, 0x33, 0x20,
	0x0C, 0x06, 0x07, 0x34, 0x3E, 0x35, 0x45, 0x5B, 0x0D, 0x5D, 0x19, 0x3C,
	0x3F, 0x71, 0x5E, 0x15, 0x45, 0x59, 0x17, 0x29, 0x26, 0x3F, 0x0D, 0x38,
	0x28, 0x0E, 0x5D, 0x3B, 0x17, 0x05, 0x2C, 0x34, 0x13, 0x7B, 0x3C, 0x2D,
	0x09, 0x39, 0x03, 0x02, 0x50, 0x2F, 0x32, 0x3A, 0x5B, 0x14, 0x00, 0x05,
	0x24, 0x0B, 0x25, 0x04, 0x09, 0x29, 0x3B, 0x2C, 0x5C, 0x11, 0x03, 0x20,
	0x2C, 0x21, 0x5C, 0x05, 0x1F, 0x58, 0x5E, 0x07, 0x12, 0x5F, 0x37, 0x0D,
	0x31, 0x75, 0x2F, 0x08, 0x29, 0x5E, 0x76, 0x20, 0x26, 0x1C, 0x52, 0x72,
	0x01, 0x52, 0x5E, 0x27, 0x05, 0x1E, 0x4A, 0x37, 0x0D, 0x16, 0x5A, 0x4E,
	0x04, 0x58, 0x10, 0x0F, 0x0F, 0x3F, 0x5E, 0x3B, 0x27, 0x08, 0x0F, 0x03,
	0x38, 0x26, 0x36, 0x21, 0x20, 0x73, 0x23, 0x09, 0x3C, 0x01, 0x0B, 0x0B,
	0x10, 0x3C, 0x05, 0x35, 0x22, 0x2C, 0x0A, 0x5E, 0x30, 0x1D, 0x02, 0x28,
	0x5C, 0x18, 0x5C, 0x39, 0x03, 0x08, 0x00, 0x1D, 0x59, 0x17, 0x5E, 0x0F,
	0x5C, 0x10, 0x3A, 0x3D, 0x01, 0x29, 0x02, 0x2A, 0x31, 0x2C, 0x01, 0x05,
	0x56, 0x5F, 0x0A, 0x19, 0x00, 0x2D, 0x2A, 0x74, 0x08, 0x50, 0x14, 0x01,
	0x23, 0x22, 0x23, 0x26, 0x2C, 0x13, 0x43, 0x17, 0x5F, 0x39, 0x0F, 0x24,
	0x2F, 0x3E, 0x5F, 0x74, 0x43, 0x11, 0x27, 0x06, 0x21, 0x08, 0x54, 0x5B,
	0x18, 0x14, 0x08, 0x53, 0x20, 0x44, 0x32, 0x2A, 0x1B, 0x0C, 0x44, 0x2A,
	0x19, 0x04, 0x41, 0x13, 0x20, 0x5A, 0x0B, 0x59, 0x3A, 0x7A, 0x05, 0x4E,
	0x01, 0x3F, 0x3A, 0x05, 0x08, 0x5A, 0x3F, 0x77, 0x22, 0x53, 0x17, 0x28,
	0x7B, 0x47, 0x11, 0x3E, 0x2F, 0x6D, 0x34, 0x14, 0x3C, 0x09, 0x0A, 0x55,
	0x27, 0x14, 0x40, 0x2B, 0x00, 0x00, 0x3B, 0x44, 0x72, 0x21, 0x10, 0x57,
	0x59, 0x0F, 0x1E, 0x4E, 0x09, 0x20, 0x13, 0x1F, 0x50, 0x38, 0x33, 0x0F,
	0x05, 0x25, 0x22, 0x3A, 0x33, 0x03, 0x2A, 0x0B, 0x2E, 0x04, 0x3B, 0x4A,
	0x5A, 0x01, 0x77, 0x3F, 0x0F, 0x0F, 0x1F, 0x2A, 0x05, 0x10, 0x1B, 0x1A,
	0x33, 0x24, 0x06, 0x29, 0x1B, 0x73, 0x59, 0x4E, 0x26, 0x26, 0x71, 0x2A,
	0x51, 0x37, 0x3A, 0x17, 0x15, 0x05, 0x0A, 0x52, 0x38, 0x0E, 0x19, 0x5E,
	0x3B, 0x1A, 0x43, 0x23, 0x5A, 0x5E, 0x6D, 0x5A, 0x11, 0x01, 0x07, 0x72,
	0x1F, 0x00, 0x0A, 0x52, 0x29, 0x5B, 0x05, 0x1B, 0x31, 0x7B, 0x1F, 0x55,
	0x58, 0x02, 0x10, 0x39, 0x2E, 0x45, 0x2F, 0x71, 0x47, 0x27, 0x05, 0x5B,
	0x72, 0x06, 0x29, 0x45, 0x1F, 0x38, 0x04, 0x59, 0x1F, 0x5E, 0x0B, 0x1B,
	0x11, 0x19, 0x3E, 0x38, 0x06, 0x20, 0x0C, 0x58, 0x27, 0x0A, 0x2F, 0x21,
	0x22, 0x24, 0x54, 0x35, 0x2F, 0x33, 0x2E, 0x01, 0x0F, 0x09, 0x1B, 0x69,
	0x08, 0x07, 0x39, 0x31, 0x0A, 0x43, 0x09, 0x1F, 0x3E, 0x03, 0x22, 0x59,
	0x0A, 0x3A, 0x0C, 0x47, 0x50, 0x0C, 0x08, 0x00, 0x09, 0x59, 0x5F, 0x3A,
	0x0D, 0x0A, 0x0C, 0x3C, 0x18, 0x74, 0x16, 0x39, 0x59, 0x1B, 0x29, 0x0B,
	0x04, 0x5C, 0x02, 0x69, 0x21, 0x07, 0x3E, 0x21, 0x70, 0x27, 0x50, 0x56,
	0x53, 0x0F, 0x1B, 0x50, 0x02, 0x07, 0x27, 0x2B, 0x07, 0x24, 0x5B, 0x23,
	0x54, 0x09, 0x5F, 0x3D, 0x20, 0x5E, 0x54, 0x07, 0x12, 0x06, 0x08, 0x07,
	0x21, 0x04, 0x32, 0x59, 0x0B, 0x5D, 0x26, 0x14, 0x02, 0x59, 0x2F, 0x1C,
	0x21, 0x28, 0x55, 0x02, 0x5F, 0x04, 0x38, 0x56, 0x20, 0x2F, 0x07, 0x2B,
	0x13, 0x3B, 0x5F, 0x75, 0x14, 0x0E, 0x2F, 0x31, 0x20, 0x0A, 0x06, 0x1D,
	0x06, 0x2D, 0x2D, 0x3B, 0x5B, 0x5D, 0x32, 0x1D, 0x30, 0x29, 0x2A, 0x3B,
	0x2E, 0x19, 0x23, 0x2C, 0x38, 0x14, 0x23, 0x01, 0x04, 0x73, 0x38, 0x07,
	0x5E, 0x3F, 0x06, 0x3D, 0x03, 0x04, 0x40, 0x28, 0x08, 0x07, 0x24, 0x2F,
	0x72, 0x23, 0x10, 0x5C, 0x18, 0x29, 0x5A, 0x08, 0x1C, 0x59, 0x14, 0x39,
	0x1B, 0x14, 0x59, 0x31, 0x36, 0x2A, 0x34, 0x0C, 0x74, 0x2B, 0x26, 0x59,
	0x0E, 0x29, 0x16, 0x37, 0x0B, 0x52, 0x28, 0x23, 0x04, 0x04, 0x0C, 0x2B,
	0x1F, 0x0E, 0x0B, 0x0D, 0x00, 0x59, 0x04, 0x3F, 0x1D, 0x16, 0x2E, 0x1B,
	0x5E, 0x20, 0x25, 0x5A, 0x29, 0x5F, 0x39, 0x06, 0x5F, 0x2D, 0x2D, 0x32,
	0x0A, 0x1F, 0x17, 0x5C, 0x20, 0x77, 0x1C, 0x2E, 0x5A, 0x11, 0x15, 0x1F,
	0x56, 0x0B, 0x38, 0x00, 0x03, 0x08, 0x58, 0x5E, 0x07, 0x0B, 0x00, 0x57,
	0x00, 0x1A, 0x1E, 0x29, 0x5A, 0x19, 0x30, 0x35, 0x4A, 0x0C, 0x3A, 0x2E,
	0x15, 0x0F, 0x20, 0x3B, 0x1A, 0x5C, 0x2E, 0x17, 0x1F, 0x0F, 0x5E, 0x0C,
	0x18, 0x05, 0x0F, 0x5A, 0x24, 0x2D, 0x2F, 0x7A, 0x47, 0x2B, 0x23, 0x39,
	0x14, 0x1F, 0x1B, 0x3E, 0x59, 0x0C, 0x2D, 0x0C, 0x00, 0x11, 0x74, 0x18,
	0x29, 0x38, 0x29, 0x10, 0x36, 0x04, 0x3F, 0x2E, 0x2F, 0x19, 0x27, 0x2D,
	0x0D, 0x13, 0x01, 0x24, 0x03, 0x31, 0x00, 0x3B, 0x37, 0x5A, 0x1D, 0x23,
	0x5A, 0x17, 0x5A, 0x01, 0x76, 0x35, 0x4E, 0x45, 0x02, 0x3B, 0x20, 0x31,
	0x1E, 0x04, 0x2A, 0x3F, 0x04, 0x3D, 0x03, 0x10, 0x5F, 0x37, 0x41, 0x3B,
	0x3A, 0x05, 0x31, 0x2D, 0x0E, 0x0C, 0x14, 0x07, 0x58, 0x3E, 0x0E, 0x19,
	0x20, 0x34, 0x3F, 0x06, 0x34, 0x2A, 0x08, 0x28, 0x13, 0x20, 0x0E, 0x27,
	0x59, 0x2E, 0x3B, 0x0B, 0x57, 0x3D, 0x76, 0x24, 0x29, 0x57, 0x52, 0x6D,
	0x3B, 0x0B, 0x1A, 0x3A, 0x10, 0x28, 0x52, 0x1A, 0x32, 0x7A, 0x27, 0x04,
	0x29, 0x07, 0x2E, 0x3C, 0x56, 0x56, 0x31, 0x1A, 0x55, 0x16, 0x3A, 0x28,
	0x74, 0x07, 0x0B, 0x28, 0x21, 0x77, 0x5E, 0x0E, 0x0F, 0x2C, 0x7A, 0x15,
	0x00, 0x04, 0x38, 0x03, 0x38, 0x4A, 0x59, 0x1F, 0x01, 0x19, 0x4E, 0x38,
	0x5E, 0x74, 0x04, 0x50, 0x0C, 0x04, 0x21, 0x43, 0x0C, 0x0D, 0x5B, 0x07,
	0x5C, 0x4A, 0x0D, 0x22, 0x2B, 0x03, 0x58, 0x3F, 0x3B, 0x13, 0x21, 0x2F,
	0x14, 0x23, 0x28, 0x09, 0x05, 0x02, 0x08, 0x12, 0x2B, 0x18, 0x5D, 0x58,
	0x12, 0x55, 0x0F, 0x0C, 0x39, 0x2D, 0x1A, 0x0F, 0x2A, 0x3C, 0x11, 0x0A,
	0x58, 0x5E, 0x40, 0x0A, 0x05, 0x09, 0x28, 0x04, 0x2D, 0x3D, 0x53, 0x0C,
	0x09, 0x72, 0x0F, 0x26, 0x2F, 0x00, 0x72, 0x0E, 0x30, 0x5C, 0x59, 0x6D,
	0x28, 0x50, 0x25, 0x2D, 0x37, 0x19, 0x19, 0x37, 0x0E, 0x0A, 0x08, 0x28,
	0x08, 0x2D, 0x35, 0x3D, 0x59, 0x0B, 0x03, 0x0E, 0x18, 0x22, 0x18, 0x06,
	0x0A, 0x29, 0x2C, 0x56, 0x28, 0x16, 0x1D, 0x30, 0x21, 0x24, 0x16, 0x54,
	0x02, 0x2F, 0x08, 0x11, 0x04, 0x52, 0x3F, 0x13, 0x72, 0x03, 0x26, 0x05,
	0x21, 0x16, 0x0A, 0x28, 0x5A, 0x3D, 0x26, 0x1D, 0x26, 0x45, 0x27, 0x2E,
	0x5E, 0x27, 0x03, 0x09, 0x73, 0x29, 0x32, 0x3F, 0x1E, 0x3A, 0x1A, 0x0F,
	0x39, 0x2D, 0x09, 0x2D, 0x0C, 0x58, 0x19, 0x38, 0x35, 0x33, 0x02, 0x39,
	0x33, 0x02, 0x2A, 0x59, 0x19, 0x13, 0x04, 0x53, 0x22, 0x22, 0x6D, 0x47,
	0x23, 0x5F, 0x0E, 0x32, 0x43, 0x2F, 0x45, 0x01, 0x0F, 0x38, 0x14, 0x5F,
	0x04, 0x33, 0x58, 0x55, 0x5C, 0x3F, 0x36, 0x1E, 0x2E, 0x5B, 0x58, 0x6D,
	0x25, 0x19, 0x14, 0x2E, 0x71, 0x02, 0x08, 0x36, 0x3C, 0x00, 0x18, 0x15,
	0x1F, 0x0A, 0x05, 0x5C, 0x32, 0x2A, 0x5C, 0x13, 0x16, 0x4E, 0x04, 0x02,
	0x2B, 0x27, 0x4A, 0x57, 0x28, 0x01, 0x43, 0x37, 0x56, 0x58, 0x15, 0x55,
	0x2F, 0x59, 0x2D, 0x23, 0x0D, 0x18, 0x25, 0x5F, 0x0C, 0x1A, 0x35, 0x37,
	0x13, 0x2F, 0x5F, 0x17, 0x3C, 0x1A, 0x35, 0x22, 0x50, 0x59, 0x2F, 0x12,
	0x3D, 0x05, 0x06, 0x26, 0x7B, 0x1C, 0x29, 0x19, 0x06, 0x18, 0x07, 0x52,
	0x01, 0x04, 0x21, 0x36, 0x39, 0x18, 0x0A, 0x07, 0x3C, 0x12, 0x23, 0x19,
	0x21, 0x35, 0x38, 0x36, 0x03, 0x70, 0x5E, 0x0D, 0x2A, 0x3F, 0x20, 0x1C,
	0x59, 0x2C, 0x3B, 0x7A, 0x16, 0x36, 0x34, 0x5A, 0x0B, 0x55, 0x28, 0x29,
	0x53, 0x33, 0x39, 0x30, 0x14, 0x07, 0x10, 0x07, 0x58, 0x38, 0x2F, 0x28,
	0x28, 0x03, 0x5D, 0x33, 0x05, 0x29, 0x34, 0x5F, 0x25, 0x2E, 0x22, 0x50,
	0x5D, 0x20, 0x2E, 0x1E, 0x10, 0x00, 0x1E, 0x2A, 0x09, 0x52, 0x36, 0x2A,
	0x0D, 0x59, 0x39, 0x0F, 0x13, 0x71, 0x29, 0x35, 0x2A, 0x0A, 0x37, 0x0E,
	0x13, 0x58, 0x2C, 0x25, 0x34, 0x15, 0x18, 0x1F, 0x72, 0x0F, 0x26, 0x1A,
	0x3B, 0x2C, 0x26, 0x2D, 0x0C, 0x07, 0x21, 0x34, 0x06, 0x17, 0x31, 0x05,
	0x06, 0x11, 0x25, 0x32, 0x23, 0x59, 0x25, 0x03, 0x0F, 0x06, 0x38, 0x33,
	0x1B, 0x32, 0x2E, 0x3E, 0x0B, 0x57, 0x22, 0x03, 0x21, 0x23, 0x02, 0x2E,
	0x7B, 0x2A, 0x0B, 0x22, 0x0E, 0x77, 0x5A, 0x2F, 0x5F, 0x19, 0x35, 0x1D,
	0x19, 0x39, 0x02, 0x36, 0x0F, 0x20, 0x3D, 0x1B, 0x6D, 0x3D, 0x24, 0x22,
	0x05, 0x70, 0x5C, 0x29, 0x24, 0x32, 0x36, 0x24, 0x1B, 0x00, 0x2F, 0x33,
	0x3D, 0x0B, 0x07, 0x5D, 0x34, 0x03, 0x06, 0x2B, 0x52, 0x17, 0x1A, 0x55,
	0x37, 0x59, 0x24, 0x1B, 0x30, 0x08, 0x1B, 0x77, 0x5A, 0x11, 0x01, 0x1F,
	0x71, 0x19, 0x57, 0x0D, 0x0E, 0x25, 0x04, 0x59, 0x01, 0x25, 0x35, 0x58,
	0x25, 0x0C, 0x01, 0x35, 0x39, 0x03, 0x36, 0x44, 0x3B, 0x0A, 0x25, 0x58,
	0x21, 0x2B, 0x28, 0x35, 0x1B, 0x12, 0x2F, 0x2F, 0x0A, 0x19, 0x13, 0x07,
	0x59, 0x0B, 0x22, 0x04, 0x21, 0x2E, 0x08, 0x1E, 0x3F, 0x70, 0x5B, 0x30,
	0x0B, 0x3C, 0x75, 0x26, 0x15, 0x39, 0x58, 0x10, 0x3E, 0x11, 0x08, 0x5D,
	0x0A, 0x15, 0x22, 0x5C, 0x5C, 0x09, 0x25, 0x20, 0x2C, 0x5D, 0x1A, 0x0E,
	0x0B, 0x5A, 0x26, 0x70, 0x38, 0x55, 0x08, 0x5E, 0x2A, 0x1A, 0x0E, 0x2B,
	0x59, 0x24, 0x3D, 0x15, 0x5D, 0x2D, 0x32, 0x2E, 0x29, 0x01, 0x26, 0x10,
	0x2F, 0x56, 0x17, 0x52, 0x10, 0x1E, 0x36, 0x0B, 0x5A, 0x30, 0x07, 0x55,
	0x19, 0x1E, 0x0E, 0x01, 0x2A, 0x27, 0x22, 0x04, 0x0A, 0x31, 0x0C, 0x21,
	0x21, 0x3B, 0x1B, 0x2B, 0x52, 0x0A, 0x0F, 0x12, 0x14, 0x01, 0x25, 0x27,
	0x0D, 0x06, 0x5E, 0x72, 0x3B, 0x11, 0x1D, 0x18, 0x0A, 0x27, 0x0D, 0x18,
	0x27, 0x07, 0x59, 0x35, 0x26, 0x19, 0x33, 0x2A, 0x30, 0x2C, 0x0D, 0x17,
	0x54, 0x0D, 0x21, 0x52, 0x76, 0x43, 0x2B, 0x41, 0x0D, 0x34, 0x58, 0x0B,
	0x17, 0x2C, 0x1A, 0x3E, 0x56, 0x56, 0x27, 0x7A, 0x27, 0x39, 0x21, 0x1E,
	0x7B, 0x0D, 0x02, 0x3B, 0x5F, 0x0E, 0x5F, 0x57, 0x5A, 0x04, 0x29, 0x1B,
	0x27, 0x00, 0x08, 0x2C, 0x55, 0x24, 0x58, 0x52, 0x70, 0x2E, 0x34, 0x3B,
	0x5B, 0x13, 0x1D, 0x07, 0x2A, 0x20, 0x26, 0x1F, 0x09, 0x5F, 0x39, 0x32,
	0x3E, 0x54, 0x2F, 0x2E, 0x38, 0x21, 0x26, 0x28, 0x0F, 0x38, 0x3E, 0x2C,
	0x1B, 0x1D, 0x09, 0x3E, 0x27, 0x3D, 0x29, 0x74, 0x3C, 0x39, 0x1F, 0x09,
	0x08, 0x29, 0x0B, 0x5F, 0x3D, 0x2B, 0x02, 0x33, 0x0F, 0x5B, 0x34, 0x1C,
	0x12, 0x2B, 0x1A, 0x70, 0x03, 0x33, 0x5C, 0x1A, 0x76, 0x14, 0x17, 0x0A,
	0x02, 0x75, 0x36, 0x18, 0x28, 0x13, 0x10, 0x0F, 0x09, 0x3F, 0x3E, 0x0E,
	0x20, 0x53, 0x3E, 0x5A, 0x27, 0x23, 0x33, 0x0D, 0x2C, 0x24, 0x00, 0x0A,
	0x21, 0x20, 0x0C, 0x14, 0x32, 0x29, 0x3E, 0x70, 0x1E, 0x2D, 0x5A, 0x52,
	0x08, 0x29, 0x10, 0x45, 0x2F, 0x2F, 0x05, 0x08, 0x07, 0x3B, 0x28, 0x3A,
	0x36, 0x05, 0x38, 0x1B, 0x2D, 0x38, 0x09, 0x1C, 0x6D, 0x16, 0x0E, 0x08,
	0x29, 0x28, 0x20, 0x54, 0x5F, 0x0C, 0x2B, 0x3D, 0x56, 0x3A, 0x40, 0x0D,
	0x15, 0x50, 0x1B, 0x06, 0x16, 0x43, 0x52, 0x05, 0x2E, 0x31, 0x25, 0x14,
	0x3B, 0x2C, 0x0A, 0x21, 0x38, 0x00, 0x1D, 0x10, 0x08, 0x34, 0x1E, 0x22,
	0x00, 0x1A, 0x03, 0x56, 0x1F, 0x00, 0x25, 0x10, 0x04, 0x2A, 0x09, 0x09,
	0x14, 0x2C, 0x5B, 0x32, 0x3B, 0x29, 0x5E, 0x08, 0x09, 0x18, 0x18, 0x21,
	0x28, 0x23, 0x5F, 0x37, 0x1B, 0x33, 0x2B, 0x2A, 0x0C, 0x5B, 0x5E, 0x33,
	0x28, 0x0D, 0x59, 0x5A, 0x3A, 0x0D, 0x15, 0x1E, 0x0E, 0x0B, 0x34, 0x03,
	0x19, 0x1A, 0x2D, 0x2A, 0x13, 0x14, 0x28, 0x10, 0x18, 0x1B, 0x01, 0x0E,
	0x30, 0x16, 0x20, 0x57, 0x1A, 0x38, 0x03, 0x00, 0x1C, 0x40, 0x0E, 0x14,
	0x57, 0x18, 0x19, 0x38, 0x03, 0x04, 0x3A, 0x3C, 0x27, 0x47, 0x12, 0x23,
	0x0E, 0x30, 0x20, 0x18, 0x04, 0x5E, 0x75, 0x28, 0x3B, 0x21, 0x3E, 0x14,
	0x00, 0x2A, 0x34, 0x08, 0x38, 0x36, 0x24, 0x1B, 0x26, 0x28, 0x34, 0x19,
	0x57, 0x09, 0x21, 0x21, 0x2D, 0x2B, 0x5A, 0x77, 0x23, 0x34, 0x1A, 0x3F,
	0x1A, 0x18, 0x28, 0x3C, 0x03, 0x2D, 0x5A, 0x17, 0x26, 0x5F, 0x1A, 0x1D,
	0x53, 0x05, 0x5D, 0x13, 0x59, 0x0A, 0x1A, 0x38, 0x34, 0x24, 0x13, 0x5D,
	0x0F, 0x7B, 0x1D, 0x00, 0x57, 0x3C, 0x31, 0x19, 0x0B, 0x24, 0x28, 0x27,
	0x14, 0x29, 0x22, 0x1D, 0x36, 0x2B, 0x08, 0x18, 0x21, 0x01, 0x59, 0x12,
	0x5A, 0x09, 0x72, 0x3C, 0x39, 0x59, 0x58, 0x21, 0x03, 0x09, 0x05, 0x12,
	0x73, 0x2A, 0x39, 0x20, 0x08, 0x0B, 0x3A, 0x07, 0x1F, 0x3A, 0x14, 0x58,
	0x09, 0x38, 0x38, 0x30, 0x3C, 0x0E, 0x20, 0x33, 0x72, 0x38, 0x35, 0x45,
	0x5E, 0x2F, 0x28, 0x31, 0x24, 0x12, 0x24, 0x34, 0x38, 0x3D, 0x59, 0x31,
	0x5A, 0x59, 0x5D, 0x3B, 0x17, 0x18, 0x05, 0x14, 0x18, 0x0D, 0x19, 0x15,
	0x19, 0x0A, 0x75, 0x34, 0x17, 0x5A, 0x00, 0x23, 0x20, 0x0F, 0x3D, 0x52,
	0x0F, 0x03, 0x04, 0x58, 0x19, 0x25, 0x28, 0x28, 0x03, 0x3D, 0x04, 0x59,
	0x2A, 0x20, 0x3A, 0x28, 0x5D, 0x07, 0x3E, 0x44, 0x36, 0x0D, 0x37, 0x5E,
	0x27, 0x21, 0x38, 0x11, 0x59, 0x5A, 0x08, 0x16, 0x0C, 0x00, 0x2D, 0x1B,
	0x06, 0x24, 0x05, 0x00, 0x2E, 0x14, 0x53, 0x2C, 0x26, 0x33, 0x55, 0x50,
	0x0F, 0x25, 0x71, 0x08, 0x08, 0x24, 0x19, 0x73, 0x36, 0x1B, 0x29, 0x18,
	0x37, 0x5F, 0x4E, 0x2A, 0x3D, 0x6D, 0x19, 0x17, 0x06, 0x19, 0x32, 0x3E,
	0x59, 0x02, 0x3C, 0x2D, 0x2B, 0x16, 0x1A, 0x5C, 0x75, 0x29, 0x3B, 0x0B,
	0x1F, 0x70, 0x59, 0x59, 0x5E, 0x03, 0x20, 0x5A, 0x2E, 0x04, 0x0D, 0x31,
	0x5A, 0x56, 0x3F, 0x0E, 0x34, 0x14, 0x56, 0x0D, 0x5C, 0x15, 0x18, 0x07,
	0x29, 0x5B, 0x30, 0x5E, 0x00, 0x27, 0x00, 0x3A, 0x21, 0x52, 0x14, 0x5E,
	0x01, 0x2E, 0x2E, 0x5A, 0x00, 0x29, 0x02, 0x0C, 0x07, 0x12, 0x6D, 0x25,
	0x10, 0x21, 0x5C, 0x69, 0x3F, 0x35, 0x05, 0x0C, 0x28, 0x0A, 0x26, 0x22,
	0x22, 0x0C, 0x47, 0x39, 0x05, 0x5A, 0x34, 0x1D, 0x0E, 0x0A, 0x08, 0x75,
	0x5E, 0x12, 0x3E, 0x22, 0x32, 0x14, 0x00, 0x08, 0x44, 0x09, 0x1F, 0x58,
	0x0C, 0x28, 0x77, 0x5F, 0x55, 0x1E, 0x3B, 0x71, 0x5E, 0x12, 0x00, 0x3D,
	0x14, 0x43, 0x52, 0x03, 0x0E, 0x04, 0x06, 0x3B, 0x1A, 0x44, 0x0A, 0x22,
	0x2A, 0x45, 0x5B, 0x10, 0x1C, 0x54, 0x18, 0x13, 0x71, 0x29, 0x52, 0x05,
	0x40, 0x15, 0x39, 0x2A, 0x3D, 0x38, 0x00, 0x1E, 0x11, 0x41, 0x01, 0x10,
	0x58, 0x58, 0x3D, 0x3C, 0x2F, 0x1D, 0x50, 0x1D, 0x20, 0x29, 0x38, 0x08,
	0x34, 0x1C, 0x7A, 0x08, 0x52, 0x05, 0x53, 0x72, 0x0B, 0x57, 0x19, 0x1F,
	0x26, 0x3E, 0x55, 0x1A, 0x5B, 0x0F, 0x5E, 0x59, 0x5B, 0x53, 0x72, 0x03,
	0x58, 0x06, 0x33, 0x04, 0x1B, 0x12, 0x2F, 0x26, 0x7A, 0x1F, 0x23, 0x5A,
	0x2F, 0x2C, 0x59, 0x27, 0x04, 0x0C, 0x07, 0x47, 0x0C, 0x5D, 0x0D, 0x31,
	0x3C, 0x19, 0x5A, 0x12, 0x05, 0x06, 0x00, 0x14, 0x13, 0x1B, 0x18, 0x27,
	0x08, 0x05, 0x04, 0x58, 0x33, 0x5C, 0x40, 0x03, 0x36, 0x16, 0x25, 0x13,
	0x2F, 0x25, 0x30, 0x1B, 0x3B, 0x0C, 0x28, 0x17, 0x3A, 0x04, 0x71, 0x00,
	0x0C, 0x24, 0x5A, 0x21, 0x58, 0x2A, 0x06, 0x1D, 0x14, 0x28, 0x08, 0x21,
	0x32, 0x69, 0x55, 0x32, 0x1A, 0x25, 0x7A, 0x5C, 0x56, 0x3A, 0x08, 0x0E,
	0x58, 0x18, 0x23, 0x53, 0x6D, 0x06, 0x33, 0x5C, 0x5D, 0x6D, 0x0D, 0x29,
	0x1D, 0x28, 0x23, 0x1C, 0x27, 0x2A, 0x1E, 0x3B, 0x28, 0x10, 0x5C, 0x59,
	0x2E, 0x23, 0x2B, 0x0B, 0x40, 0x27, 0x58, 0x11, 0x06, 0x2E, 0x07, 0x5D,
	0x2E, 0x5E, 0x3B, 0x69, 0x26, 0x23, 0x0A, 0x40, 0x2A, 0x1E, 0x18, 0x5E,
	0x3B, 0x2A, 0x05, 0x00, 0x3C, 0x2F, 0x7B, 0x28, 0x35, 0x06, 0x58, 0x71,
	0x01, 0x10, 0x0C, 0x1C, 0x74, 0x2D, 0x4A, 0x5B, 0x25, 0x2C, 0x3B, 0x33,
	0x28, 0x1B, 0x2A, 0x04, 0x29, 0x01, 0x1D, 0x21, 0x54, 0x2F, 0x0A, 0x5D,
	0x26, 0x1E, 0x14, 0x2D, 0x07, 0x16, 0x03, 0x34, 0x3A, 0x5B, 0x24, 0x20,
	0x08, 0x56, 0x24, 0x69, 0x14, 0x53, 0x2C, 0x2D, 0x0C, 0x19, 0x0A, 0x3A,
	0x02, 0x2E, 0x3B, 0x0A, 0x3C, 0x02, 0x24, 0x06, 0x53, 0x36, 0x3C, 0x25,
	0x0A, 0x17, 0x3F, 0x23, 0x04, 0x5A, 0x36, 0x18, 0x29, 0x05, 0x07, 0x4E,
	0x41, 0x58, 0x34, 0x03, 0x19, 0x5F, 0x03, 0x24, 0x2D, 0x56, 0x1E, 0x5B,
	0x05, 0x5A, 0x50, 0x3D, 0x03, 0x11, 0x2E, 0x31, 0x20, 0x38, 0x05, 0x0B,
	0x12, 0x03, 0x12, 0x11, 0x58, 0x0D, 0x0D, 0x38, 0x17, 0x23, 0x2C, 0x05,
	0x5B, 0x17, 0x06, 0x56, 0x2D, 0x25, 0x30, 0x54, 0x03, 0x1E, 0x5F, 0x10,
	0x1B, 0x26, 0x3D, 0x5D, 0x12, 0x2D, 0x59, 0x2A, 0x0F, 0x2B, 0x38, 0x38,
	0x18, 0x26, 0x2E, 0x34, 0x55, 0x0D, 0x04, 0x2F, 0x34, 0x03, 0x3A, 0x11,
	0x31, 0x5F, 0x05, 0x0C, 0x3D, 0x75, 0x08, 0x22, 0x27, 0x08, 0x12, 0x15,
	0x36, 0x25, 0x18, 0x7A, 0x23, 0x58, 0x0C, 0x1A, 0x14, 0x5E, 0x31, 0x1A,
	0x07, 0x32, 0x5D, 0x59, 0x17, 0x31, 0x0E, 0x2E, 0x51, 0x24, 0x19, 0x16,
	0x06, 0x51, 0x19, 0x33, 0x06, 0x15, 0x34, 0x37, 0x1E, 0x01, 0x1C, 0x39,
	0x07, 0x5E, 0x2E, 0x5F, 0x03, 0x56, 0x25, 0x73, 0x15, 0x2C, 0x0B, 0x5E,
	0x26, 0x0B, 0x38, 0x05, 0x44, 0x6D, 0x5A, 0x35, 0x5E, 0x07, 0x26, 0x34,
	0x17, 0x16, 0x20, 0x21, 0x28, 0x59, 0x3F, 0x20, 0x71, 0x0B, 0x26, 0x2D,
	0x09, 0x06, 0x14, 0x20, 0x0D, 0x2E, 0x74, 0x1A, 0x22, 0x0B, 0x38, 0x14,
	0x1C, 0x58, 0x14, 0x3A, 0x1B, 0x1E, 0x2C, 0x01, 0x12, 0x72, 0x5A, 0x09,
	0x59, 0x38, 0x14, 0x1E, 0x29, 0x05, 0x32, 0x32, 0x09, 0x52, 0x5B, 0x18,
	0x7B, 0x06, 0x16, 0x23, 0x0D, 0x24, 0x2D, 0x23, 0x09, 0x32, 0x04, 0x3C,
	0x4E, 0x27, 0x3F, 0x03, 0x03, 0x0E, 0x20, 0x29, 0x18, 0x05, 0x24, 0x0C,
	0x5B, 0x0D, 0x2D, 0x0A, 0x2F, 0x21, 0x35, 0x1E, 0x26, 0x2F, 0x1C, 0x0C,
	0x01, 0x4A, 0x20, 0x04, 0x77, 0x05, 0x0E, 0x18, 0x0D, 0x14, 0x05, 0x51,
	0x04, 0x08, 0x14, 0x5C, 0x2A, 0x22, 0x01, 0x0D, 0x58, 0x37, 0x17, 0x09,
	0x33, 0x04, 0x0B, 0x37, 0x00, 0x27, 0x38, 0x08, 0x34, 0x52, 0x03, 0x22,
	0x52, 0x0C, 0x20, 0x20, 0x20, 0x52, 0x05, 0x28, 0x0E, 0x1D, 0x03, 0x16,
	0x2C, 0x77, 0x3C, 0x08, 0x3C, 0x2D, 0x21, 0x00, 0x3B, 0x17, 0x59, 0x27,
	0x2B, 0x52, 0x2C, 0x32, 0x14, 0x1D, 0x3B, 0x03, 0x53, 0x27, 0x59, 0x56,
	0x39, 0x29, 0x32, 0x03, 0x2F, 0x59, 0x38, 0x36, 0x27, 0x13, 0x09, 0x12,
	0x7B, 0x22, 0x09, 0x0C, 0x5C, 0x0D, 0x1F, 0x3B, 0x58, 0x2C, 0x12, 0x15,
	0x53, 0x1C, 0x05, 0x17, 0x5D, 0x4A, 0x2B, 0x09, 0x77, 0x01, 0x2B, 0x08,
	0x25, 0x70, 0x04, 0x58, 0x08, 0x31, 0x34, 0x5A, 0x10, 0x1D, 0x5E, 0x00,
	0x08, 0x1B, 0x08, 0x1D, 0x77, 0x2B, 0x2B, 0x37, 0x31, 0x20, 0x14, 0x0B,
	0x0A, 0x53, 0x74, 0x00, 0x08, 0x2F, 0x1A, 0x2E, 0x04, 0x59, 0x25, 0x05,
	0x6D, 0x3C, 0x3B, 0x3E, 0x53, 0x01, 0x01, 0x26, 0x0F, 0x0E, 0x0E, 0x03,
	0x29, 0x27, 0x31, 0x2C, 0x2B, 0x0E, 0x1B, 0x27, 0x2E, 0x24, 0x2D, 0x2F,
	0x3A, 0x0B, 0x55, 0x39, 0x0F, 0x21, 0x2B, 0x1B, 0x06, 0x2B, 0x58, 0x7B,
	0x03, 0x52, 0x2B, 0x18, 0x3B, 0x21, 0x20, 0x07, 0x03, 0x2A, 0x0B, 0x03,
	0x18, 0x06, 0x08, 0x1A, 0x36, 0x0F, 0x38, 0x31, 0x47, 0x27, 0x23, 0x32,
	0x36, 0x27, 0x22, 0x34, 0x00, 0x08, 0x1C, 0x3B, 0x3C, 0x3A, 0x05, 0x3A,
	0x24, 0x2A, 0x26, 0x2D, 0x0D, 0x06, 0x07, 0x06, 0x0E, 0x21, 0x20, 0x5C,
	0x2A, 0x17, 0x1F, 0x30, 0x0D, 0x58, 0x09, 0x0F, 0x3B, 0x45, 0x2F, 0x06,
	0x18, 0x38, 0x04, 0x23, 0x24, 0x5C, 0x54, 0x09, 0x52, 0x2E, 0x3E, 0x23,
	0x07, 0x5B, 0x14, 0x3E, 0x2A, 0x3B, 0x1A, 0x14, 0x05, 0x23, 0x19, 0x19,
	0x0E, 0x02, 0x50, 0x27, 0x26, 0x18, 0x39, 0x18, 0x3F, 0x31, 0x1B, 0x47,
	0x13, 0x5B, 0x3A, 0x36, 0x28, 0x06, 0x3D, 0x5B, 0x0F, 0x2E, 0x18, 0x16,
	0x2C, 0x2C, 0x3A, 0x06, 0x2D, 0x2A, 0x76, 0x1E, 0x0F, 0x04, 0x28, 0x34,
	0x36, 0x2C, 0x2B, 0x12, 0x01, 0x28, 0x54, 0x18, 0x0A, 0x2F, 0x3F, 0x03,
	0x25, 0x59, 0x2B, 0x3E, 0x2F, 0x1E, 0x2F, 0x35, 0x00, 0x2F, 0x1A, 0x44,
	0x2B, 0x1C, 0x25, 0x27, 0x38, 0x77, 0x5D, 0x29, 0x24, 0x5D, 0x3B, 0x0B,
	0x30, 0x22, 0x06, 0x3B, 0x59, 0x35, 0x0A, 0x04, 0x71, 0x5D, 0x4A, 0x34,
	0x1E, 0x25, 0x2F, 0x51, 0x23, 0x32, 0x01, 0x54, 0x20, 0x45, 0x3F, 0x73,
	0x26, 0x37, 0x23, 0x19, 0x20, 0x27, 0x31, 0x16, 0x5D, 0x18, 0x23, 0x11,
	0x07, 0x5D, 0x38, 0x3F, 0x24, 0x39, 0x0A, 0x2E, 0x55, 0x22, 0x58, 0x27,
	0x26, 0x34, 0x06, 0x00, 0x32, 0x28, 0x3D, 0x20, 0x17, 0x58, 0x21, 0x1E,
	0x54, 0x5F, 0x04, 0x36, 0x23, 0x16, 0x1C, 0x1D, 0x38, 0x3D, 0x1B, 0x05,
	0x24, 0x0F, 0x55, 0x13, 0x41, 0x0C, 0x06, 0x23, 0x13, 0x19, 0x38, 0x37,
	0x21, 0x02, 0x3C, 0x38, 0x29, 0x25, 0x04, 0x38, 0x5F, 0x05, 0x59, 0x54,
	0x1E, 0x1A, 0x69, 0x26, 0x19, 0x41, 0x5A, 0x03, 0x3B, 0x04, 0x2C, 0x2E,
	0x3B, 0x47, 0x56, 0x56, 0x2C, 0x1B, 0x27, 0x24, 0x1B, 0x40, 0x26, 0x14,
	0x07, 0x0C, 0x27, 0x2B, 0x03, 0x17, 0x27, 0x09, 0x30, 0x36, 0x00, 0x25,
	0x44, 0x0F, 0x07, 0x16, 0x59, 0x58, 0x10, 0x21, 0x18, 0x0A, 0x21, 0x10,
	0x39, 0x22, 0x5C, 0x5F, 0x20, 0x27, 0x0A, 0x22, 0x11, 0x01, 0x5B, 0x0E,
	0x3C, 0x52, 0x13, 0x01, 0x02, 0x1C, 0x52, 0x3B, 0x3C, 0x53, 0x29, 0x02,
	0x0B, 0x43, 0x11, 0x34, 0x1F, 0x09, 0x2D, 0x12, 0x2A, 0x31, 0x77, 0x1E,
	0x23, 0x5F, 0x38, 0x05, 0x06, 0x16, 0x18, 0x20, 0x2D, 0x26, 0x52, 0x56,
	0x40, 0x35, 0x38, 0x0F, 0x36, 0x19, 0x36, 0x5C, 0x38, 0x0D, 0x18, 0x33,
	0x24, 0x25, 0x0B, 0x05, 0x09, 0x04, 0x05, 0x45, 0x2F, 0x24, 0x22, 0x12,
	0x3F, 0x5E, 0x24, 0x0F, 0x25, 0x0D, 0x39, 0x2F, 0x21, 0x29, 0x01, 0x21,
	0x35, 0x0B, 0x17, 0x04, 0x5B, 0x01, 0x2B, 0x23, 0x0D, 0x07, 0x21, 0x2E,
	0x00, 0x2B, 0x32, 0x07, 0x09, 0x02, 0x39, 0x11, 0x33, 0x29, 0x29, 0x0C,
	0x5B, 0x2B, 0x55, 0x16, 0x28, 0x0F, 0x03, 0x54, 0x17, 0x45, 0x5F, 0x0D,
	0x1D, 0x27, 0x57, 0x0F, 0x03, 0x34, 0x4E, 0x39, 0x5F, 0x6D, 0x08, 0x00,
	0x0B, 0x0E, 0x75, 0x35, 0x2F, 0x3C, 0x3D, 0x32, 0x02, 0x57, 0x45, 0x29,
	0x38, 0x47, 0x0C, 0x59, 0x27, 0x29, 0x2E, 0x30, 0x20, 0x31, 0x36, 0x5D,
	0x0B, 0x01, 0x5B, 0x24, 0x5E, 0x22, 0x59, 0x04, 0x16, 0x34, 0x08, 0x19,
	0x02, 0x01, 0x1B, 0x52, 0x5F, 0x08, 0x30, 0x3B, 0x11, 0x5D, 0x29, 0x70,
	0x1A, 0x53, 0x38, 0x1C, 0x14, 0x47, 0x18, 0x41, 0x21, 0x25, 0x14, 0x20,
	0x41, 0x2A, 0x07, 0x3A, 0x1B, 0x00, 0x1D, 0x75, 0x5E, 0x31, 0x1B, 0x25,
	0x27, 0x20, 0x59, 0x37, 0x5F, 0x77, 0x0D, 0x2C, 0x3A, 0x32, 0x0F, 0x0E,
	0x15, 0x07, 0x3F, 0x2D, 0x2B, 0x22, 0x0B, 0x09, 0x0F, 0x0B, 0x4A, 0x2B,
	0x04, 0x18, 0x05, 0x26, 0x05, 0x24, 0x2A, 0x05, 0x2A, 0x26, 0x08, 0x05,
	0x5E, 0x2E, 0x03, 0x07, 0x16, 0x01, 0x1B, 0x05, 0x0C, 0x23, 0x0A, 0x30,
	0x18, 0x1F, 0x2D, 0x2F, 0x56, 0x39, 0x2A, 0x28, 0x28, 0x00, 0x56, 0x0A,
	0x06, 0x2F, 0x32, 0x24, 0x38, 0x0A, 0x5B, 0x0E, 0x14, 0x18, 0x6D, 0x26,
	0x20, 0x00, 0x32, 0x1B, 0x3E, 0x3B, 0x5B, 0x18, 0x12, 0x27, 0x16, 0x03,
	0x06, 0x76, 0x58, 0x25, 0x00, 0x07, 0x18, 0x21, 0x2F, 0x38, 0x2C, 0x7B,
	0x0D, 0x37, 0x3C, 0x1D, 0x09, 0x47, 0x23, 0x5C, 0x3B, 0x38, 0x16, 0x25,
	0x27, 0x59, 0x72, 0x0B, 0x39, 0x06, 0x18, 0x21, 0x19, 0x2C, 0x3C, 0x02,
	0x0F, 0x3A, 0x36, 0x17, 0x59, 0x04, 0x1C, 0x51, 0x2C, 0x06, 0x20, 0x02,
	0x0B, 0x3C, 0x1B, 0x74, 0x21, 0x52, 0x3A, 0x5A, 0x6D, 0x1C, 0x12, 0x1A,
	0x2D, 0x36, 0x1D, 0x57, 0x01, 0x25, 0x16, 0x24, 0x38, 0x5D, 0x24, 0x36,
	0x0E, 0x2F, 0x3B, 0x38, 0x32, 0x09, 0x59, 0x2B, 0x20, 0x13, 0x22, 0x36,
	0x00, 0x40, 0x21, 0x23, 0x38, 0x03, 0x3C, 0x0E, 0x35, 0x11, 0x38, 0x11,
	0x26, 0x15, 0x25, 0x59, 0x58, 0x3A, 0x0D, 0x19, 0x02, 0x01, 0x2B, 0x07,
	0x06, 0x21, 0x02, 0x7A, 0x38, 0x2B, 0x58, 0x3F, 0x05, 0x55, 0x23, 0x04,
	0x13, 0x14, 0x34, 0x4A, 0x2B, 0x1C, 0x2D, 0x19, 0x38, 0x21, 0x26, 0x04,
	0x3E, 0x39, 0x3A, 0x1E, 0x14, 0x1D, 0x11, 0x45, 0x03, 0x37, 0x03, 0x0A,
	0x09, 0x5A, 0x2D, 0x00, 0x0E, 0x5F, 0x12, 0x3B, 0x04, 0x16, 0x2B, 0x0D,
	0x73, 0x36, 0x0C, 0x5E, 0x13, 0x31, 0x43, 0x19, 0x3E, 0x5C, 0x2A, 0x0F,
	0x13, 0x24, 0x3D, 0x03, 0x34, 0x2D, 0x19, 0x52, 0x72, 0x3B, 0x22, 0x3F,
	0x1B, 0x35, 0x0A, 0x30, 0x0D, 0x21, 0x2C, 0x39, 0x11, 0x58, 0x03, 0x36,
	0x3C, 0x14, 0x45, 0x40, 0x01, 0x2B, 0x51, 0x3B, 0x1F, 0x1B, 0x5F, 0x0F,
	0x5D, 0x3E, 0x2D, 0x39, 0x08, 0x1B, 0x02, 0x03, 0x0D, 0x4A, 0x0B, 0x02,
	0x01, 0x20, 0x24, 0x19, 0x20, 0x29, 0x01, 0x53, 0x38, 0x09, 0x2D, 0x2D,
	0x51, 0x07, 0x22, 0x13, 0x07, 0x23, 0x00, 0x32, 0x2F, 0x05, 0x28, 0x41,
	0x12, 0x2D, 0x36, 0x28, 0x5D, 0x0F, 0x11, 0x5A, 0x2D, 0x3B, 0x03, 0x1A,
	0x03, 0x30, 0x19, 0x04, 0x09, 0x58, 0x22, 0x2D, 0x52, 0x3A, 0x0E, 0x0C,
	0x5B, 0x05, 0x25, 0x2F, 0x4A, 0x0C, 0x24, 0x31, 0x00, 0x12, 0x1D, 0x1D,
	0x28, 0x0E, 0x2B, 0x14, 0x11, 0x14, 0x36, 0x2D, 0x45, 0x08, 0x2D, 0x3B,
	0x56, 0x26, 0x3B, 0x69, 0x35, 0x57, 0x2B, 0x40, 0x74, 0x5B, 0x50, 0x2B,
	0x1E, 0x21, 0x28, 0x32, 0x16, 0x09, 0x37, 0x08, 0x08, 0x0B, 0x0C, 0x10,
	0x0A, 0x18, 0x38, 0x44, 0x25, 0x21, 0x2F, 0x34, 0x5F, 0x15, 0x2F, 0x32,
	0x58, 0x0F, 0x28, 0x5D, 0x06, 0x2C, 0x0D, 0x6D, 0x1C, 0x0E, 0x36, 0x20,
	0x77, 0x06, 0x36, 0x20, 0x1D, 0x0F, 0x47, 0x28, 0x23, 0x39, 0x28, 0x15,
	0x34, 0x19, 0x39, 0x34, 0x0F, 0x0F, 0x45, 0x5F, 0x0E, 0x19, 0x35, 0x3C,
	0x2C, 0x75, 0x3D, 0x07, 0x57, 0x00, 0x7B, 0x3D, 0x0F, 0x09, 0x31, 0x05,
	0x58, 0x26, 0x00, 0x24, 0x0A, 0x5D, 0x2A, 0x37, 0x05, 0x0D, 0x21, 0x54,
	0x00, 0x31, 0x7B, 0x2D, 0x25, 0x58, 0x5B, 0x2D, 0x0E, 0x11, 0x16, 0x3E,
	0x77, 0x18, 0x23, 0x24, 0x0E, 0x30, 0x05, 0x29, 0x45, 0x0A, 0x75, 0x3D,
	0x38, 0x1B, 0x04, 0x2D, 0x04, 0x54, 0x57, 0x2C, 0x05, 0x54, 0x51, 0x00,
	0x3D, 0x06, 0x0A, 0x2E, 0x2B, 0x1D, 0x23, 0x29, 0x38, 0x2A, 0x5B, 0x32,
	0x2B, 0x09, 0x0B, 0x26, 0x3B, 0x47, 0x09, 0x22, 0x25, 0x7B, 0x05, 0x2B,
	0x45, 0x23, 0x0D, 0x2E, 0x56, 0x34, 0x3A, 0x2D, 0x5B, 0x57, 0x5D, 0x2F,
	0x34, 0x19, 0x57, 0x2F, 0x3A, 0x2D, 0x34, 0x58, 0x59, 0x31, 0x2C, 0x5D,
	0x2F, 0x1B, 0x07, 0x36, 0x47, 0x15, 0x04, 0x1A, 0x23, 0x19, 0x38, 0x5E,
	0x33, 0x70, 0x36, 0x52, 0x0A, 0x05, 0x6D, 0x2B, 0x4A, 0x59, 0x3B, 0x3A,
	0x5A, 0x1B, 0x0B, 0x33, 0x07, 0x58, 0x10, 0x04, 0x0D, 0x08, 0x1B, 0x25,
	0x02, 0x20, 0x04, 0x16, 0x07, 0x1A, 0x5F, 0x38, 0x2D, 0x33, 0x5F, 0x0D,
	0x3A, 0x5A, 0x57, 0x45, 0x2D, 0x3B, 0x21, 0x30, 0x24, 0x38, 0x69, 0x55,
	0x50, 0x5E, 0x0C, 0x25, 0x14, 0x2A, 0x36, 0x2A, 0x00, 0x05, 0x25, 0x28,
	0x2C, 0x0B, 0x3B, 0x18, 0x59, 0x3D, 0x29, 0x28, 0x36, 0x1E, 0x20, 0x3B,
	0x34, 0x22, 0x5D, 0x39, 0x24, 0x25, 0x0A, 0x08, 0x1B, 0x29, 0x2A, 0x10,
	0x0D, 0x1B, 0x70, 0x27, 0x23, 0x00, 0x2E, 0x36, 0x2F, 0x14, 0x5F, 0x0A,
	0x17, 0x0F, 0x20, 0x56, 0x0C, 0x00, 0x0F, 0x22, 0x09, 0x03, 0x21, 0x54,
	0x06, 0x3B, 0x5A, 0x17, 0x5C, 0x2F, 0x5B, 0x26, 0x28, 0x21, 0x29, 0x38,
	0x2C, 0x14, 0x5C, 0x55, 0x2B, 0x25, 0x2E, 0x36, 0x27, 0x1F, 0x06, 0x73,
	0x2A, 0x54, 0x36, 0x1B, 0x13, 0x21, 0x23, 0x5A, 0x2F, 0x34, 0x21, 0x2A,
	0x59, 0x5C, 0x1B, 0x01, 0x24, 0x2F, 0x0C, 0x75, 0x5B, 0x10, 0x28, 0x2C,
	0x2F, 0x47, 0x27, 0x00, 0x06, 0x2F, 0x16, 0x2C, 0x16, 0x1D, 0x30, 0x34,
	0x04, 0x0F, 0x22, 0x35, 0x1C, 0x11, 0x0C, 0x12, 0x2B, 0x59, 0x4E, 0x3D,
	0x1E, 0x13, 0x3C, 0x52, 0x37, 0x05, 0x08, 0x25, 0x2E, 0x19, 0x3F, 0x28,
	0x18, 0x0A, 0x00, 0x0D, 0x25, 0x1E, 0x32, 0x03, 0x32, 0x04, 0x25, 0x13,
	0x3F, 0x2A, 0x12, 0x09, 0x07, 0x36, 0x26, 0x6D, 0x25, 0x0A, 0x57, 0x5E,
	0x21, 0x19, 0x2B, 0x0B, 0x25, 0x0F, 0x2A, 0x30, 0x19, 0x2E, 0x36, 0x29,
	0x25, 0x38, 0x59, 0x15, 0x47, 0x15, 0x20, 0x40, 0x25, 0x23, 0x14, 0x20,
	0x2E, 0x75, 0x58, 0x31, 0x05, 0x11, 0x73, 0x5F, 0x05, 0x22, 0x20, 0x77,
	0x15, 0x20, 0x59, 0x20, 0x18, 0x1F, 0x17, 0x16, 0x1A, 0x71, 0x23, 0x52,
	0x06, 0x31, 0x1A, 0x3B, 0x17, 0x1A, 0x32, 0x6D, 0x3F, 0x38, 0x20, 0x06,
	0x0C, 0x5E, 0x04, 0x3C, 0x04, 0x0B, 0x1C, 0x4E, 0x3E, 0x12, 0x24, 0x23,
	0x17, 0x39, 0x18, 0x2A, 0x1D, 0x09, 0x45, 0x3F, 0x28, 0x0A, 0x12, 0x04,
	0x08, 0x06, 0x54, 0x2C, 0x1E, 0x3F, 0x23, 0x2E, 0x2A, 0x03, 0x2E, 0x0D,
	0x26, 0x16, 0x2A, 0x29, 0x71, 0x14, 0x22, 0x1A, 0x27, 0x73, 0x25, 0x10,
	0x5F, 0x5D, 0x2C, 0x36, 0x52, 0x38, 0x5B, 0x09, 0x04, 0x56, 0x04, 0x1E,
	0x37, 0x08, 0x18, 0x06, 0x12, 0x7A, 0x47, 0x4E, 0x19, 0x3A, 0x0F, 0x2A,
	0x56, 0x1A, 0x39, 0x6D, 0x58, 0x52, 0x16, 0x22, 0x32, 0x54, 0x0B, 0x3B,
	0x5D, 0x21, 0x2D, 0x2F, 0x22, 0x21, 0x10, 0x20, 0x34, 0x2D, 0x09, 0x7B,
	0x5E, 0x2C, 0x07, 0x5D, 0x2B, 0x21, 0x14, 0x23, 0x5F, 0x03, 0x3E, 0x06,
	0x21, 0x40, 0x16, 0x58, 0x18, 0x0C, 0x29, 0x31, 0x23, 0x54, 0x16, 0x18,
	0x05, 0x39, 0x2A, 0x3F, 0x0E, 0x15, 0x3F, 0x0A, 0x22, 0x02, 0x74, 0x5C,
	0x57, 0x07, 0x02, 0x75, 0x2A, 0x15, 0x2F, 0x39, 0x0D, 0x0D, 0x14, 0x5D,
	0x2F, 0x7B, 0x1B, 0x14, 0x1D, 0x23, 0x32, 0x02, 0x26, 0x20, 0x23, 0x7B,
	0x29, 0x02, 0x0A, 0x33, 0x76, 0x07, 0x35, 0x23, 0x12, 0x74, 0x15, 0x53,
	0x34, 0x5E, 0x74, 0x5E, 0x3B, 0x5F, 0x5E, 0x32, 0x2B, 0x0A, 0x36, 0x19,
	0x29, 0x09, 0x08, 0x1D, 0x2A, 0x0F, 0x27, 0x2C, 0x2F, 0x18, 0x0A, 0x2A,
	0x57, 0x18, 0x21, 0x38, 0x14, 0x34, 0x02, 0x52, 0x30, 0x27, 0x55, 0x25,
	0x11, 0x2F, 0x0D, 0x54, 0x2C, 0x22, 0x11, 0x20, 0x15, 0x29, 0x2F, 0x08,
	0x38, 0x50, 0x5F, 0x3A, 0x21, 0x2A, 0x23, 0x19, 0x04, 0x33, 0x1F, 0x0A,
	0x28, 0x2D, 0x7A, 0x2E, 0x38, 0x14, 0x25, 0x74, 0x24, 0x37, 0x29, 0x13,
	0x25, 0x01, 0x18, 0x22, 0x38, 0x34, 0x28, 0x0C, 0x19, 0x18, 0x32, 0x07,
	0x0A, 0x2B, 0x28, 0x10, 0x55, 0x15, 0x3F, 0x3C, 0x18, 0x1F, 0x12, 0x14,
	0x32, 0x14, 0x39, 0x57, 0x5B, 0x2C, 0x33, 0x22, 0x36, 0x34, 0x5F, 0x3B,
	0x39, 0x1B, 0x0F, 0x24, 0x04, 0x23, 0x37, 0x28, 0x23, 0x12, 0x1E, 0x02,
	0x1E, 0x01, 0x27, 0x27, 0x05, 0x26, 0x3F, 0x38, 0x59, 0x56, 0x07, 0x1C,
	0x0D, 0x5F, 0x05, 0x03, 0x40, 0x29, 0x3F, 0x14, 0x5D, 0x3A, 0x77, 0x22,
	0x26, 0x1B, 0x11, 0x04, 0x3F, 0x04, 0x06, 0x0D, 0x3A, 0x27, 0x27, 0x41,
	0x5B, 0x1A, 0x07, 0x13, 0x1A, 0x1C, 0x7A, 0x58, 0x4E, 0x16, 0x20, 0x30,
	0x0D, 0x16, 0x0D, 0x58, 0x1A, 0x0F, 0x56, 0x3E, 0x28, 0x0C, 0x0B, 0x12,
	0x3A, 0x5F, 0x0B, 0x1B, 0x34, 0x18, 0x22, 0x7A, 0x1F, 0x29, 0x22, 0x39,
	0x37, 0x39, 0x2E, 0x3B, 0x01, 0x18, 0x34, 0x04, 0x2C, 0x2C, 0x69, 0x5E,
	0x24, 0x38, 0x29, 0x73, 0x2D, 0x30, 0x5B, 0x23, 0x24, 0x3F, 0x22, 0x09,
	0x02, 0x24, 0x55, 0x36, 0x5F, 0x40, 0x74, 0x2D, 0x02, 0x04, 0x24, 0x3A,
	0x5F, 0x19, 0x5D, 0x1A, 0x31, 0x3D, 0x55, 0x05, 0x25, 0x14, 0x3C, 0x33,
	0x26, 0x26, 0x09, 0x55, 0x0F, 0x56, 0x53, 0x08, 0x58, 0x37, 0x59, 0x21,
	0x10, 0x3E, 0x03, 0x5B, 0x5A, 0x12, 0x0F, 0x27, 0x37, 0x29, 0x18, 0x3D,
	0x37, 0x22, 0x05, 0x30, 0x38, 0x25, 0x3A, 0x1D, 0x0E, 0x03, 0x0E, 0x03,
	0x03, 0x04, 0x3F, 0x04, 0x34, 0x2A, 0x25, 0x1C, 0x16, 0x37, 0x38, 0x2D,
	0x08, 0x2F, 0x5A, 0x2F, 0x27, 0x20, 0x37, 0x2F, 0x1D, 0x31, 0x2B, 0x22,
	0x0A, 0x24, 0x38, 0x3F, 0x09, 0x16, 0x01, 0x6D, 0x05, 0x13, 0x07, 0x08,
	0x17, 0x14, 0x05, 0x2B, 0x5E, 0x25, 0x3C, 0x09, 0x2F, 0x38, 0x13, 0x0F,
	0x12, 0x1B, 0x00, 0x0E, 0x3B, 0x09, 0x56, 0x24, 0x15, 0x3D, 0x2F, 0x24,
	0x31, 0x0A, 0x02, 0x54, 0x0F, 0x12, 0x1B, 0x1D, 0x27, 0x03, 0x0F, 0x2A,
	0x2A, 0x03, 0x03, 0x31, 0x69, 0x36, 0x56, 0x41, 0x21, 0x00, 0x5B, 0x2D,
	0x2A, 0x12, 0x69, 0x0A, 0x03, 0x3F, 0x39, 0x09, 0x1E, 0x28, 0x3D, 0x44,
	0x2E, 0x1F, 0x17, 0x3F, 0x2E, 0x04, 0x26, 0x0F, 0x17, 0x31, 0x7B, 0x1B,
	0x33, 0x38, 0x1E, 0x21, 0x0D, 0x09, 0x0C, 0x03, 0x21, 0x5E, 0x2B, 0x58,
	0x1E, 0x0F, 0x1B, 0x09, 0x0A, 0x02, 0x2C, 0x43, 0x05, 0x3F, 0x20, 0x0A,
	0x36, 0x28, 0x1D, 0x0C, 0x17, 0x24, 0x24, 0x45, 0x00, 0x2F, 0x3A, 0x4A,
	0x1F, 0x01, 0x2F, 0x21, 0x31, 0x36, 0x19, 0x18, 0x1B, 0x0C, 0x2B, 0x2F,
	0x69, 0x00, 0x32, 0x0B, 0x0D, 0x2A, 0x2E, 0x03, 0x0B, 0x21, 0x31, 0x1B,
	0x36, 0x3B, 0x25, 0x31, 0x3A, 0x53, 0x0D, 0x3E, 0x1A, 0x55, 0x28, 0x2D,
	0x20, 0x2C, 0x24, 0x33, 0x16, 0x24, 0x15, 0x54, 0x54, 0x16, 0x1E, 0x7A,
	0x47, 0x22, 0x39, 0x33, 0x38, 0x5F, 0x17, 0x21, 0x5B, 0x04, 0x34, 0x34,
	0x37, 0x5C, 0x3B, 0x02, 0x29, 0x18, 0x08, 0x76, 0x1D, 0x11, 0x3B, 0x44,
	0x6D, 0x0B, 0x11, 0x36, 0x18, 0x7A, 0x25, 0x23, 0x1D, 0x1B, 0x72, 0x14,
	0x57, 0x21, 0x02, 0x31, 0x1C, 0x25, 0x5A, 0x2D, 0x03, 0x5F, 0x26, 0x26,
	0x29, 0x0D, 0x5D, 0x20, 0x1C, 0x3E, 0x33, 0x2A, 0x27, 0x59, 0x59, 0x0F,
	0x54, 0x4E, 0x56, 0x24, 0x18, 0x3B, 0x57, 0x2D, 0x03, 0x34, 0x24, 0x0A,
	0x0C, 0x09, 0x2D, 0x2F, 0x18, 0x23, 0x0A, 0x73, 0x5E, 0x31, 0x07, 0x25,
	0x35, 0x14, 0x2B, 0x1D, 0x3C, 0x21, 0x21, 0x26, 0x56, 0x39, 0x74, 0x5C,
	0x12, 0x25, 0x22, 0x25, 0x25, 0x37, 0x04, 0x59, 0x04, 0x3F, 0x0B, 0x27,
	0x5D, 0x30, 0x2B, 0x07, 0x09, 0x2C, 0x24, 0x3D, 0x37, 0x39, 0x3F, 0x28,
	0x09, 0x23, 0x25, 0x5F, 0x1B, 0x04, 0x56, 0x5E, 0x11, 0x14, 0x3F, 0x37,
	0x37, 0x1C, 0x35, 0x15, 0x02, 0x5D, 0x59, 0x31, 0x3D, 0x11, 0x2D, 0x28,
	0x76, 0x43, 0x59, 0x26, 0x33, 0x37, 0x21, 0x29, 0x45, 0x25, 0x73, 0x00,
	0x4E, 0x21, 0x04, 0x24, 0x38, 0x55, 0x3D, 0x29, 0x35, 0x08, 0x51, 0x25,
	0x0A, 0x38, 0x5C, 0x18, 0x29, 0x2F, 0x0C, 0x5C, 0x39, 0x34, 0x5F, 0x0C,
	0x27, 0x4A, 0x56, 0x3D, 0x18, 0x29, 0x19, 0x26, 0x23, 0x36, 0x29, 0x55,
	0x34, 0x5E, 0x36, 0x5E, 0x00, 0x1A, 0x58, 0x77, 0x27, 0x50, 0x16, 0x53,
	0x20, 0x16, 0x2E, 0x01, 0x3D, 0x75, 0x1F, 0x16, 0x21, 0x18, 0x35, 0x2D,
	0x4E, 0x1E, 0x33, 0x71, 0x47, 0x08, 0x21, 0x0D, 0x33, 0x35, 0x34, 0x21,
	0x40, 0x10, 0x19, 0x2F, 0x01, 0x1E, 0x20, 0x14, 0x26, 0x2C, 0x0D, 0x0E,
	0x26, 0x59, 0x0C, 0x2D, 0x01, 0x05, 0x54, 0x41, 0x0C, 0x2F, 0x06, 0x3B,
	0x39, 0x0F, 0x03, 0x1F, 0x50, 0x0C, 0x0C, 0x23, 0x20, 0x0D, 0x07, 0x07,
	0x72, 0x1D, 0x0D, 0x17, 0x33, 0x01, 0x1B, 0x57, 0x1A, 0x38, 0x7A, 0x2B,
	0x2D, 0x24, 0x2A, 0x0D, 0x1C, 0x2B, 0x08, 0x09, 0x77, 0x2B, 0x02, 0x2A,
	0x3D, 0x2E, 0x08, 0x0F, 0x14, 0x3B, 0x0B, 0x0E, 0x54, 0x5D, 0x03, 0x34,
	0x38, 0x33, 0x2D, 0x5E, 0x36, 0x06, 0x0F, 0x3D, 0x19, 0x26, 0x08, 0x3B,
	0x1E, 0x3E, 0x23, 0x1E, 0x57, 0x5C, 0x38, 0x0E, 0x06, 0x00, 0x1B, 0x13,
	0x21, 0x0A, 0x14, 0x17, 0x02, 0x7A, 0x5B, 0x51, 0x2F, 0x3D, 0x77, 0x23,
	0x2E, 0x45, 0x26, 0x73, 0x21, 0x19, 0x2F, 0x1A, 0x06, 0x19, 0x04, 0x45,
	0x5D, 0x21, 0x34, 0x25, 0x06, 0x1F, 0x28, 0x07, 0x39, 0x23, 0x5F, 0x2F,
	0x3C, 0x16, 0x04, 0x2E, 0x14, 0x21, 0x14, 0x36, 0x2F, 0x0D, 0x1A, 0x24,
	0x22, 0x0A, 0x38, 0x0D, 0x29, 0x29, 0x08, 0x7B, 0x2A, 0x24, 0x02, 0x20,
	0x2F, 0x2A, 0x57, 0x0D, 0x25, 0x00, 0x20, 0x04, 0x3C, 0x53, 0x0A, 0x5B,
	0x2A, 0x26, 0x19, 0x24, 0x5C, 0x05, 0x26, 0x3F, 0x69, 0x5E, 0x09, 0x5A,
	0x23, 0x72, 0x5F, 0x17, 0x04, 0x44, 0x16, 0x58, 0x52, 0x09, 0x01, 0x34,
	0x06, 0x07, 0x3C, 0x40, 0x15, 0x58, 0x4E, 0x18, 0x3F, 0x24, 0x28, 0x04,
	0x3C, 0x24, 0x6D, 0x0A, 0x25, 0x1C, 0x5E, 0x71, 0x47, 0x36, 0x24, 0x08,
	0x6D, 0x1C, 0x09, 0x09, 0x20, 0x17, 0x1F, 0x11, 0x36, 0x5C, 0x0B, 0x27,
	0x2D, 0x36, 0x07, 0x34, 0x5E, 0x0D, 0x28, 0x1B, 0x07, 0x36, 0x19, 0x45,
	0x3C, 0x75, 0x2B, 0x19, 0x04, 0x5C, 0x33, 0x58, 0x06, 0x19, 0x23, 0x75,
	0x5C, 0x55, 0x1B, 0x26, 0x2B, 0x47, 0x3B, 0x25, 0x07, 0x77, 0x3B, 0x07,
	0x14, 0x52, 0x21, 0x2F, 0x23, 0x21, 0x02, 0x25, 0x0E, 0x08, 0x00, 0x3C,
	0x03, 0x1B, 0x33, 0x5A, 0x25, 0x15, 0x0D, 0x03, 0x07, 0x5E, 0x09, 0x15,
	0x2E, 0x2A, 0x52, 0x21, 0x5D, 0x10, 0x5D, 0x2E, 0x29, 0x02, 0x15, 0x37,
	0x12, 0x18, 0x19, 0x33, 0x28, 0x27, 0x20, 0x21, 0x30, 0x02, 0x27, 0x1B,
	0x2E, 0x0F, 0x41, 0x3D, 0x01, 0x55, 0x20, 0x25, 0x19, 0x06, 0x27, 0x55,
	0x1E, 0x3F, 0x07, 0x3C, 0x34, 0x24, 0x05, 0x70, 0x22, 0x2F, 0x2C, 0x39,
	0x05, 0x14, 0x08, 0x09, 0x2E, 0x28, 0x5E, 0x07, 0x0C, 0x3C, 0x71, 0x21,
	0x16, 0x17, 0x1A, 0x03, 0x43, 0x53, 0x3D, 0x03, 0x18, 0x3D, 0x32, 0x04,
	0x3D, 0x0F, 0x2E, 0x08, 0x04, 0x21, 0x31, 0x08, 0x08, 0x24, 0x5E, 0x75,
	0x14, 0x59, 0x23, 0x18, 0x2E, 0x3E, 0x2E, 0x0A, 0x5C, 0x27, 0x14, 0x2D,
	0x1E, 0x2F, 0x38, 0x54, 0x02, 0x3D, 0x21, 0x2E, 0x16, 0x52, 0x09, 0x26,
	0x76, 0x08, 0x2E, 0x0D, 0x2F, 0x73, 0x23, 0x0D, 0x09, 0x07, 0x3B, 0x01,
	0x13, 0x3D, 0x40, 0x1B, 0x00, 0x2B, 0x08, 0x3C, 0x2E, 0x54, 0x13, 0x01,
	0x09, 0x2B, 0x1A, 0x31, 0x58, 0x5A, 0x2F, 0x0D, 0x2B, 0x26, 0x22, 0x70,
	0x2E, 0x17, 0x02, 0x1A, 0x2F, 0x1B, 0x52, 0x1E, 0x2F, 0x17, 0x47, 0x15,
	0x34, 0x5F, 0x0C, 0x54, 0x00, 0x5B, 0x3B, 0x28, 0x03, 0x13, 0x2B, 0x3A,
	0x7B, 0x5C, 0x23, 0x27, 0x2D, 0x2F, 0x24, 0x50, 0x21, 0x05, 0x16, 0x04,
	0x18, 0x5D, 0x07, 0x0F, 0x23, 0x0E, 0x16, 0x02, 0x3A, 0x2B, 0x19, 0x39,
	0x3F, 0x6D, 0x59, 0x0E, 0x16, 0x2C, 0x0D, 0x24, 0x58, 0x2D, 0x59, 0x28,
	0x2D, 0x17, 0x16, 0x5F, 0x3A, 0x43, 0x53, 0x27, 0x5F, 0x71, 0x1E, 0x19,
	0x1A, 0x5A, 0x2E, 0x58, 0x31, 0x1B, 0x2A, 0x77, 0x2E, 0x35, 0x2B, 0x32,
	0x24, 0x14, 0x0E, 0x08, 0x53, 0x37, 0x25, 0x14, 0x5B, 0x0F, 0x07, 0x2A,
	0x08, 0x2B, 0x31, 0x2E, 0x28, 0x11, 0x27, 0x01, 0x1B, 0x0E, 0x50, 0x38,
	0x33, 0x2E, 0x19, 0x25, 0x1F, 0x40, 0x2C, 0x07, 0x05, 0x5C, 0x08, 0x11,
	0x3E, 0x50, 0x1D, 0x58, 0x29, 0x16, 0x0B, 0x0F, 0x20, 0x2D, 0x3E, 0x22,
	0x00, 0x2E, 0x71, 0x1D, 0x2B, 0x2D, 0x09, 0x2F, 0x06, 0x2A, 0x29, 0x39,
	0x28, 0x5D, 0x10, 0x2F, 0x28, 0x2C, 0x09, 0x15, 0x1E, 0x1A, 0x0E, 0x03,
	0x00, 0x16, 0x38, 0x36, 0x24, 0x36, 0x26, 0x1A, 0x2B, 0x3D, 0x2C, 0x2B,
	0x11, 0x07, 0x5E, 0x12, 0x58, 0x33, 0x14, 0x3C, 0x0C, 0x18, 0x39, 0x2D,
	0x0E, 0x53, 0x56, 0x53, 0x04, 0x2D, 0x09, 0x3B, 0x3E, 0x01, 0x5D, 0x29,
	0x26, 0x59, 0x12, 0x5B, 0x33, 0x39, 0x3D, 0x72, 0x3A, 0x31, 0x03, 0x3A,
	0x03, 0x5A, 0x2C, 0x45, 0x5F, 0x70, 0x0F, 0x18, 0x45, 0x5A, 0x17, 0x5A,
	0x07, 0x56, 0x27, 0x29, 0x2D, 0x27, 0x17, 0x0D, 0x7B, 0x00, 0x25, 0x19,
	0x5A, 0x13, 0x5F, 0x51, 0x19, 0x04, 0x33, 0x3A, 0x27, 0x01, 0x07, 0x03,
	0x23, 0x08, 0x57, 0x1D, 0x28, 0x5E, 0x03, 0x22, 0x25, 0x17, 0x36, 0x36,
	0x09, 0x22, 0x2C, 0x27, 0x23, 0x06, 0x3E, 0x20, 0x2A, 0x34, 0x3D, 0x05,
	0x11, 0x25, 0x13, 0x07, 0x5D, 0x05, 0x0A, 0x06, 0x5F, 0x5C, 0x2D, 0x59,
	0x08, 0x07, 0x04, 0x73, 0x06, 0x07, 0x01, 0x28, 0x37, 0x43, 0x32, 0x2C,
	0x21, 0x36, 0x35, 0x19, 0x26, 0x11, 0x71, 0x39, 0x29, 0x1E, 0x00, 0x15,
	0x47, 0x30, 0x2B, 0x1F, 0x2D, 0x0F, 0x13, 0x3F, 0x18, 0x21, 0x3D, 0x26,
	0x0D, 0x03, 0x29, 0x5F, 0x56, 0x2C, 0x44, 0x04, 0x5E, 0x23, 0x5D, 0x3F,
	0x06, 0x2D, 0x59, 0x28, 0x00, 0x31, 0x0A, 0x2F, 0x20, 0x13, 0x32, 0x2D,
	0x53, 0x3E, 0x04, 0x01, 0x3E, 0x16, 0x5D, 0x2D, 0x34, 0x05, 0x23, 0x09,
	0x0C, 0x31, 0x06, 0x0A, 0x37, 0x1C, 0x32, 0x28, 0x27, 0x3A, 0x2C, 0x12,
	0x34, 0x03, 0x3C, 0x3C, 0x0A, 0x5F, 0x28, 0x5A, 0x20, 0x38, 0x34, 0x2F,
	0x56, 0x20, 0x0B, 0x3F, 0x58, 0x3F, 0x19, 0x3B, 0x18, 0x0E, 0x24, 0x32,
	0x28, 0x26, 0x1B, 0x3D, 0x2E, 0x21, 0x39, 0x2C, 0x5B, 0x13, 0x31, 0x55,
	0x56, 0x3E, 0x0F, 0x73, 0x28, 0x55, 0x22, 0x52, 0x26, 0x19, 0x18, 0x14,
	0x5F, 0x08, 0x1B, 0x12, 0x5A, 0x22, 0x6D, 0x5F, 0x05, 0x02, 0x2E, 0x72,
	0x21, 0x17, 0x38, 0x1A, 0x11, 0x26, 0x30, 0x03, 0x0D, 0x01, 0x1F, 0x25,
	0x59, 0x00, 0x26, 0x5B, 0x2B, 0x5D, 0x2F, 0x35, 0x3F, 0x10, 0x1B, 0x19,
	0x01, 0x14, 0x25, 0x1C, 0x2E, 0x36, 0x07, 0x09, 0x22, 0x0C, 0x2A, 0x0F,
	0x0D, 0x5B, 0x33, 0x70, 0x1B, 0x03, 0x0F, 0x12, 0x2B, 0x2F, 0x10, 0x5C,
	0x3D, 0x09, 0x24, 0x11, 0x21, 0x19, 0x13, 0x16, 0x3B, 0x5A, 0x06, 0x37,
	0x0F, 0x06, 0x59, 0x0E, 0x2B, 0x1C, 0x2B, 0x16, 0x3B, 0x0C, 0x58, 0x2D,
	0x01, 0x1A, 0x17, 0x0F, 0x50, 0x2D, 0x03, 0x34, 0x16, 0x24, 0x14, 0x5E,
	0x73, 0x01, 0x00, 0x2A, 0x3D, 0x28, 0x0E, 0x2D, 0x34, 0x06, 0x2E, 0x0D,
	0x15, 0x0D, 0x52, 0x16, 0x1A, 0x59, 0x1E, 0x2E, 0x2C, 0x5A, 0x2E, 0x29,
	0x0A, 0x11, 0x00, 0x56, 0x25, 0x3E, 0x1B, 0x43, 0x13, 0x22, 0x39, 0x0E,
	0x54, 0x2B, 0x45, 0x22, 0x14, 0x06, 0x03, 0x05, 0x3E, 0x21, 0x14, 0x30,
	0x28, 0x23, 0x76, 0x24, 0x0A, 0x22, 0x2C, 0x3A, 0x38, 0x07, 0x05, 0x31,
	0x26, 0x08, 0x55, 0x18, 0x38, 0x2C, 0x19, 0x03, 0x08, 0x02, 0x0F, 0x2F,
	0x05, 0x41, 0x38, 0x24, 0x06, 0x03, 0x34, 0x0A, 0x28, 0x1A, 0x29, 0x17,
	0x1E, 0x74, 0x3D, 0x36, 0x21, 0x0A, 0x13, 0x38, 0x26, 0x2C, 0x5A, 0x07,
	0x21, 0x15, 0x5A, 0x31, 0x11, 0x2B, 0x54, 0x58, 0x28, 0x06, 0x05, 0x15,
	0x26, 0x5B, 0x2C, 0x2E, 0x2C, 0x5A, 0x07, 0x76, 0x54, 0x31, 0x2C, 0x1A,
	0x27, 0x2E, 0x2D, 0x37, 0x5C, 0x7A, 0x5E, 0x20, 0x08, 0x5C, 0x0A, 0x27,
	0x31, 0x25, 0x1A, 0x2D, 0x06, 0x22, 0x0C, 0x5E, 0x28, 0x55, 0x30, 0x1E,
	0x1D, 0x69, 0x27, 0x20, 0x34, 0x5E, 0x2F, 0x5D, 0x3B, 0x20, 0x1F, 0x00,
	0x58, 0x2B, 0x27, 0x06, 0x34, 0x3F, 0x27, 0x5F, 0x3B, 0x30, 0x22, 0x28,
	0x5A, 0x23, 0x10, 0x04, 0x03, 0x26, 0x38, 0x21, 0x1E, 0x07, 0x0C, 0x5C,
	0x15, 0x22, 0x22, 0x26, 0x09, 0x0B, 0x1E, 0x39, 0x17, 0x02, 0x3A, 0x3F,
	0x11, 0x36, 0x13, 0x2B, 0x2B, 0x09, 0x1F, 0x1C, 0x04, 0x1E, 0x20, 0x5B,
	0x1C, 0x74, 0x28, 0x12, 0x17, 0x01, 0x08, 0x02, 0x37, 0x19, 0x29, 0x00,
	0x43, 0x02, 0x1A, 0x09, 0x03, 0x0B, 0x26, 0x1B, 0x23, 0x28, 0x1E, 0x57,
	0x3B, 0x1A, 0x31, 0x47, 0x15, 0x05, 0x58, 0x71, 0x04, 0x38, 0x41, 0x1F,
	0x03, 0x03, 0x54, 0x20, 0x0F, 0x37, 0x18, 0x0B, 0x3B, 0x11, 0x0C, 0x14,
	0x57, 0x3B, 0x08, 0x14, 0x34, 0x27, 0x02, 0x44, 0x2C, 0x15, 0x38, 0x2B,
	0x20, 0x0F, 0x08, 0x02, 0x03, 0x00, 0x74, 0x29, 0x58, 0x1F, 0x09, 0x2A,
	0x55, 0x35, 0x1B, 0x5B, 0x38, 0x0E, 0x52, 0x23, 0x0A, 0x2E, 0x06, 0x18,
	0x0A, 0x53, 0x0D, 0x08, 0x38, 0x01, 0x21, 0x2E, 0x25, 0x13, 0x21, 0x0E,
	0x18, 0x21, 0x13, 0x3E, 0x53, 0x05, 0x5D, 0x39, 0x25, 0x24, 0x38, 0x38,
	0x53, 0x23, 0x3A, 0x3B, 0x07, 0x31, 0x39, 0x32, 0x7B, 0x0E, 0x23, 0x16,
	0x05, 0x32, 0x29, 0x3B, 0x2F, 0x2C, 0x00, 0x2E, 0x34, 0x37, 0x3B, 0x00,
	0x3F, 0x04, 0x1E, 0x08, 0x23, 0x3C, 0x04, 0x01, 0x2E, 0x0C, 0x2E, 0x57,
	0x0B, 0x59, 0x1A, 0x3A, 0x32, 0x0A, 0x3C, 0x04, 0x3C, 0x0C, 0x02, 0x38,
	0x13, 0x22, 0x52, 0x41, 0x09, 0x11, 0x2F, 0x06, 0x21, 0x24, 0x0A, 0x00,
	0x54, 0x5C, 0x39, 0x06, 0x0A, 0x13, 0x23, 0x27, 0x6D, 0x3D, 0x00, 0x1B,
	0x1F, 0x1A, 0x08, 0x3B, 0x1F, 0x58, 0x37, 0x16, 0x05, 0x14, 0x58, 0x15,
	0x1B, 0x32, 0x27, 0x02, 0x26, 0x04, 0x2C, 0x1F, 0x26, 0x21, 0x1C, 0x16,
	0x0A, 0x32, 0x16, 0x26, 0x57, 0x5C, 0x12, 0x20, 0x03, 0x32, 0x0B, 0x3F,
	0x04, 0x54, 0x03, 0x2A, 0x52, 0x0E, 0x3C, 0x03, 0x57, 0x5A, 0x28, 0x2E,
	0x55, 0x36, 0x18, 0x13, 0x2D, 0x07, 0x41, 0x25, 0x35, 0x03, 0x28, 0x04,
	0x44, 0x26, 0x3C, 0x0B, 0x3E, 0x25, 0x00, 0x25, 0x02, 0x28, 0x2D, 0x15,
	0x24, 0x12, 0x36, 0x1C, 0x07, 0x26, 0x11, 0x26, 0x1B, 0x77, 0x09, 0x27,
	0x28, 0x07, 0x1A, 0x0D, 0x54, 0x1B, 0x0C, 0x70, 0x19, 0x4A, 0x16, 0x5C,
	0x13, 0x0A, 0x56, 0x5B, 0x1E, 0x08, 0x08, 0x33, 0x5D, 0x2D, 0x27, 0x00,
	0x32, 0x0B, 0x2C, 0x2D, 0x03, 0x4A, 0x1E, 0x0A, 0x14, 0x3B, 0x57, 0x01,
	0x0E, 0x36, 0x23, 0x17, 0x5C, 0x1B, 0x05, 0x3B, 0x36, 0x3B, 0x39, 0x3B,
	0x0E, 0x03, 0x07, 0x13, 0x1A, 0x3E, 0x26, 0x2A, 0x12, 0x33, 0x15, 0x2A,
	0x29, 0x2D, 0x10, 0x05, 0x00, 0x28, 0x28, 0x3A, 0x07, 0x38, 0x23, 0x12,
	0x10, 0x1B, 0x54, 0x25, 0x59, 0x00, 0x5C, 0x00, 0x04, 0x3B, 0x09, 0x5B,
	0x16, 0x3F, 0x0A, 0x06, 0x0E, 0x06, 0x14, 0x3D, 0x07, 0x2E, 0x2B, 0x2A,
	0x38, 0x15, 0x1A, 0x06, 0x0B, 0x53, 0x6D, 0x2D, 0x52, 0x06, 0x0A, 0x0A,
	0x54, 0x35, 0x57, 0x07, 0x72, 0x38, 0x50, 0x0F, 0x38, 0x04, 0x2A, 0x57,
	0x07, 0x52, 0x2B, 0x35, 0x06, 0x29, 0x33, 0x1B, 0x22, 0x50, 0x23, 0x3F,
	0x23, 0x3C, 0x58, 0x0C, 0x1D, 0x24, 0x07, 0x2A, 0x06, 0x31, 0x33, 0x55,
	0x17, 0x5B, 0x27, 0x04, 0x43, 0x30, 0x5D, 0x24, 0x17, 0x38, 0x35, 0x5E,
	0x3E, 0x2E, 0x1C, 0x2D, 0x19, 0x52, 0x05, 0x1B, 0x0F, 0x5A, 0x5A, 0x0A,
	0x2B, 0x02, 0x06, 0x1A, 0x1A, 0x3E, 0x17, 0x2D, 0x53, 0x26, 0x0B, 0x30,
	0x04, 0x1E, 0x37, 0x5D, 0x56, 0x1C, 0x1E, 0x0F, 0x34, 0x31, 0x02, 0x20,
	0x18, 0x02, 0x2F, 0x3E, 0x22, 0x0C, 0x5D, 0x02, 0x5E, 0x39, 0x36, 0x05,
	0x52, 0x20, 0x2E, 0x15, 0x22, 0x27, 0x21, 0x2E, 0x35, 0x09, 0x4E, 0x2A,
	0x02, 0x25, 0x06, 0x55, 0x59, 0x3C, 0x34, 0x1C, 0x24, 0x3D, 0x06, 0x01,
	0x5C, 0x18, 0x45, 0x09, 0x23, 0x1A, 0x50, 0x3B, 0x5F, 0x32, 0x21, 0x16,
	0x41, 0x2E, 0x09, 0x3D, 0x10, 0x01, 0x59, 0x26, 0x3F, 0x23, 0x1B, 0x31,
	0x7B, 0x3E, 0x30, 0x41, 0x23, 0x0C, 0x05, 0x54, 0x45, 0x07, 0x1B, 0x1E,
	0x19, 0x1D, 0x00, 0x0B, 0x3B, 0x19, 0x2F, 0x52, 0x2F, 0x3B, 0x18, 0x1E,
	0x52, 0x12, 0x15, 0x52, 0x2C, 0x33, 0x06, 0x05, 0x25, 0x0C, 0x31, 0x0D,
	0x07, 0x57, 0x37, 0x22, 0x74, 0x16, 0x30, 0x0F, 0x3E, 0x07, 0x24, 0x51,
	0x0B, 0x1B, 0x3A, 0x35, 0x34, 0x2D, 0x3D, 0x2D, 0x29, 0x26, 0x16, 0x1B,
	0x06, 0x03, 0x22, 0x37, 0x3B, 0x17, 0x3A, 0x25, 0x07, 0x28, 0x35, 0x5B,
	0x36, 0x05, 0x25, 0x23, 0x00, 0x03, 0x28, 0x1B, 0x15, 0x24, 0x24, 0x28,
	0x27, 0x26, 0x29, 0x52, 0x23, 0x44, 0x1A, 0x1A, 0x19, 0x3F, 0x0D, 0x08,
	0x21, 0x17, 0x17, 0x2F, 0x01, 0x55, 0x37, 0x0F, 0x0D, 0x23, 0x29, 0x10,
	0x03, 0x0F, 0x37, 0x27, 0x54, 0x56, 0x22, 0x05, 0x29, 0x2E, 0x41, 0x52,
	0x26, 0x14, 0x05, 0x1B, 0x24, 0x30, 0x28, 0x0E, 0x03, 0x19, 0x25, 0x1D,
	0x38, 0x3C, 0x5A, 0x0C, 0x27, 0x36, 0x57, 0x25, 0x77, 0x38, 0x07, 0x29,
	0x58, 0x17, 0x5E, 0x36, 0x14, 0x20, 0x36, 0x08, 0x51, 0x09, 0x2C, 0x20,
	0x59, 0x37, 0x1A, 0x0E, 0x6D, 0x04, 0x34, 0x34, 0x27, 0x77, 0x1F, 0x2B,
	0x3E, 0x0D, 0x07, 0x25, 0x36, 0x20, 0x31, 0x12, 0x58, 0x12, 0x37, 0x33,
	0x31, 0x55, 0x0D, 0x17, 0x2A, 0x07, 0x23, 0x03, 0x57, 0x01, 0x03, 0x25,
	0x0B, 0x1E, 0x09, 0x28, 0x19, 0x23, 0x5C, 0x3D, 0x18, 0x36, 0x2F, 0x0F,
	0x28, 0x30, 0x35, 0x2B, 0x14, 0x00, 0x7B, 0x25, 0x27, 0x56, 0x25, 0x14,
	0x2B, 0x0F, 0x1B, 0x2F, 0x73, 0x04, 0x50, 0x5B, 0x44, 0x30, 0x22, 0x55,
	0x26, 0x2E, 0x00, 0x36, 0x07, 0x06, 0x52, 0x09, 0x01, 0x30, 0x1F, 0x1F,
	0x3B, 0x14, 0x39, 0x27, 0x2F, 0x28, 0x18, 0x39, 0x01, 0x31, 0x13, 0x59,
	0x25, 0x1A, 0x38, 0x74, 0x08, 0x09, 0x06, 0x5A, 0x05, 0x3D, 0x20, 0x1E,
	0x40, 0x72, 0x03, 0x54, 0x58, 0x26, 0x70, 0x0E, 0x2A, 0x0B, 0x21, 0x15,
	0x5F, 0x36, 0x34, 0x38, 0x14, 0x22, 0x59, 0x3D, 0x19, 0x30, 0x0D, 0x22,
	0x06, 0x0C, 0x0C, 0x0D, 0x35, 0x05, 0x26, 0x0A, 0x5E, 0x38, 0x38, 0x06,
	0x17, 0x59, 0x09, 0x25, 0x5B, 0x08, 0x5B, 0x54, 0x05, 0x01, 0x2D, 0x0D,
	0x58, 0x59, 0x0E, 0x29, 0x3C, 0x4E, 0x1B, 0x3D, 0x2F, 0x26, 0x14, 0x16,
	0x19, 0x38, 0x34, 0x10, 0x25, 0x12, 0x70, 0x29, 0x2D, 0x1B, 0x04, 0x1A,
	0x34, 0x32, 0x3A, 0x01, 0x18, 0x0B, 0x00, 0x19, 0x53, 0x26, 0x36, 0x56,
	0x3D, 0x08, 0x10, 0x5D, 0x0A, 0x2F, 0x24, 0x69, 0x58, 0x10, 0x25, 0x3C,
	0x0F, 0x1B, 0x19, 0x1F, 0x58, 0x28, 0x0F, 0x58, 0x2B, 0x40, 0x30, 0x5B,
	0x11, 0x0C, 0x5A, 0x2A, 0x3A, 0x07, 0x34, 0x1E, 0x13, 0x5C, 0x4E, 0x03,
	0x52, 0x26, 0x08, 0x2D, 0x27, 0x52, 0x03, 0x1D, 0x57, 0x03, 0x1B, 0x34,
	0x1A, 0x24, 0x0C, 0x5D, 0x0E, 0x25, 0x28, 0x1D, 0x44, 0x73, 0x01, 0x2F,
	0x5F, 0x3C, 0x70, 0x25, 0x55, 0x2A, 0x33, 0x33, 0x19, 0x0F, 0x37, 0x3E,
	0x0B, 0x22, 0x35, 0x3E, 0x19, 0x33, 0x27, 0x59, 0x5C, 0x0E, 0x3B, 0x3D,
	0x37, 0x25, 0x3E, 0x36, 0x28, 0x59, 0x38, 0x2C, 0x00, 0x06, 0x14, 0x41,
	0x18, 0x25, 0x22, 0x0B, 0x28, 0x5D, 0x06, 0x36, 0x54, 0x3D, 0x20, 0x13,
	0x06, 0x2D, 0x27, 0x39, 0x75, 0x00, 0x35, 0x5D, 0x0E, 0x16, 0x38, 0x37,
	0x38, 0x2E, 0x31, 0x24, 0x2C, 0x00, 0x5B, 0x25, 0x1B, 0x2A, 0x07, 0x44,
	0x03, 0x09, 0x54, 0x25, 0x53, 0x13, 0x34, 0x39, 0x23, 0x5C, 0x71, 0x59,
	0x29, 0x2D, 0x1C, 0x26, 0x1C, 0x12, 0x1D, 0x08, 0x18, 0x55, 0x25, 0x3D,
	0x31, 0x13, 0x2D, 0x4E, 0x09, 0x29, 0x31, 0x1A, 0x57, 0x07, 0x33, 0x7B,
	0x00, 0x2E, 0x29, 0x27, 0x2D, 0x3C, 0x20, 0x03, 0x08, 0x28, 0x1F, 0x25,
	0x1E, 0x21, 0x0F, 0x1B, 0x10, 0x1B, 0x5A, 0x73, 0x1C, 0x56, 0x1A, 0x22,
	0x6D, 0x21, 0x1B, 0x2D, 0x2C, 0x0E, 0x08, 0x2F, 0x3C, 0x52, 0x26, 0x24,
	0x4E, 0x09, 0x0E, 0x24, 0x55, 0x1B, 0x36, 0x0C, 0x77, 0x5A, 0x2B, 0x3B,
	0x27, 0x24, 0x06, 0x37, 0x1B, 0x25, 0x17, 0x02, 0x20, 0x01, 0x2D, 0x2D,
	0x5A, 0x31, 0x5B, 0x24, 0x35, 0x08, 0x59, 0x37, 0x2A, 0x69, 0x25, 0x20,
	0x22, 0x26, 0x37, 0x01, 0x33, 0x3C, 0x12, 0x05, 0x36, 0x00, 0x5D, 0x28,
	0x01, 0x28, 0x26, 0x2D, 0x2D, 0x3A, 0x03, 0x51, 0x5F, 0x0C, 0x28, 0x54,
	0x29, 0x58, 0x1A, 0x15, 0x59, 0x12, 0x2B, 0x19, 0x70, 0x35, 0x25, 0x24,
	0x2C, 0x0D, 0x05, 0x3B, 0x09, 0x44, 0x69, 0x28, 0x03, 0x5C, 0x00, 0x70,
	0x3C, 0x23, 0x21, 0x5E, 0x76, 0x28, 0x2F, 0x37, 0x26, 0x25, 0x1F, 0x0C,
	0x19, 0x5D, 0x12, 0x00, 0x0E, 0x39, 0x22, 0x25, 0x38, 0x34, 0x28, 0x3B,
	0x10, 0x5E, 0x13, 0x5F, 0x5B, 0x17, 0x0A, 0x58, 0x3B, 0x08, 0x09, 0x1D,
	0x38, 0x08, 0x2D, 0x13, 0x3E, 0x07, 0x02, 0x3D, 0x06, 0x25, 0x55, 0x0A,
	0x1D, 0x0C, 0x0A, 0x03, 0x16, 0x3A, 0x18, 0x3C, 0x30, 0x3B, 0x59, 0x71,
	0x04, 0x0C, 0x1E, 0x1A, 0x09, 0x1F, 0x39, 0x57, 0x22, 0x2C, 0x5E, 0x17,
	0x2D, 0x24, 0x01, 0x2F, 0x28, 0x1A, 0x04, 0x27, 0x0F, 0x39, 0x39, 0x27,
	0x25, 0x0F, 0x2B, 0x00, 0x5C, 0x30, 0x21, 0x37, 0x14, 0x5B, 0x75, 0x04,
	0x52, 0x41, 0x2F, 0x2E, 0x23, 0x2A, 0x18, 0x52, 0x06, 0x3F, 0x03, 0x3C,
	0x0D, 0x7A, 0x20, 0x0A, 0x07, 0x22, 0x75, 0x24, 0x4E, 0x04, 0x1A, 0x29,
	0x5A, 0x04, 0x0C, 0x02, 0x74, 0x39, 0x2E, 0x02, 0x3E, 0x29, 0x2B, 0x00,
	0x00, 0x3C, 0x06, 0x5D, 0x08, 0x07, 0x06, 0x2B, 0x5D, 0x54, 0x1C, 0x0C,
	0x33, 0x0F, 0x57, 0x3E, 0x0F, 0x2C, 0x2D, 0x06, 0x28, 0x31, 0x10, 0x02,
	0x50, 0x04, 0x1E, 0x7A, 0x03, 0x51, 0x5C, 0x5F, 0x74, 0x15, 0x27, 0x20,
	0x3F, 0x3A, 0x3C, 0x59, 0x14, 0x3E, 0x23, 0x03, 0x0A, 0x0D, 0x08, 0x23,
	0x47, 0x04, 0x02, 0x23, 0x10, 0x08, 0x04, 0x5C, 0x22, 0x75, 0x58, 0x54,
	0x3C, 0x2C, 0x2D, 0x0A, 0x15, 0x41, 0x39, 0x04, 0x3D, 0x04, 0x01, 0x2F,
	0x15, 0x01, 0x35, 0x0A, 0x1F, 0x14, 0x36, 0x0C, 0x34, 0x01, 0x27, 0x38,
	0x54, 0x29, 0x1B, 0x1A, 0x3E, 0x2A, 0x41, 0x5C, 0x0A, 0x2E, 0x00, 0x2B,
	0x24, 0x28, 0x25, 0x24, 0x59, 0x58, 0x11, 0x16, 0x2C, 0x2C, 0x00, 0x75,
	0x18, 0x37, 0x19, 0x3E, 0x77, 0x23, 0x0F, 0x34, 0x1E, 0x03, 0x1F, 0x0D,
	0x38, 0x2E, 0x77, 0x0A, 0x38, 0x2D, 0x2F, 0x2A, 0x0E, 0x0F, 0x01, 0x59,
	0x6D, 0x21, 0x15, 0x5F, 0x52, 0x06, 0x39, 0x22, 0x2A, 0x11, 0x18, 0x5D,
	0x28, 0x37, 0x21, 0x14, 0x38, 0x12, 0x57, 0x02, 0x07, 0x5E, 0x15, 0x37,
	0x20, 0x07, 0x5E, 0x4E, 0x04, 0x06, 0x73, 0x5B, 0x14, 0x5D, 0x0A, 0x29,
	0x5A, 0x35, 0x5B, 0x06, 0x06, 0x2F, 0x55, 0x21, 0x5C, 0x70, 0x14, 0x30,
	0x09, 0x2C, 0x27, 0x0E, 0x2F, 0x17, 0x2C, 0x72, 0x5A, 0x2D, 0x09, 0x1E,
	0x0A, 0x0E, 0x15, 0x28, 0x31, 0x71, 0x5F, 0x27, 0x2D, 0x23, 0x12, 0x34,
	0x25, 0x45, 0x39, 0x2E, 0x43, 0x59, 0x02, 0x04, 0x21, 0x34, 0x58, 0x2A,
	0x00, 0x3A, 0x0A, 0x19, 0x34, 0x19, 0x0D, 0x2E, 0x59, 0x07, 0x26, 0x7A,
	0x05, 0x0A, 0x24, 0x2C, 0x08, 0x0F, 0x56, 0x2F, 0x20, 0x2F, 0x04, 0x14,
	0x21, 0x5F, 0x35, 0x3F, 0x24, 0x37, 0x0D, 0x71, 0x35, 0x27, 0x16, 0x20,
	0x35, 0x3A, 0x2F, 0x08, 0x26, 0x03, 0x2B, 0x25, 0x5E, 0x18, 0x27, 0x5E,
	0x38, 0x0D, 0x0F, 0x20, 0x2E, 0x31, 0x05, 0x25, 0x13, 0x59, 0x30, 0x0B,
	0x09, 0x76, 0x26, 0x31, 0x20, 0x24, 0x2B, 0x47, 0x10, 0x57, 0x44, 0x0C,
	0x07, 0x08, 0x0F, 0x0F, 0x76, 0x16, 0x02, 0x45, 0x26, 0x0C, 0x3E, 0x50,
	0x5E, 0x1A, 0x35, 0x0D, 0x32, 0x25, 0x1C, 0x0B, 0x06, 0x19, 0x57, 0x3C,
	0x2A, 0x0E, 0x53, 0x5B, 0x1F, 0x04, 0x2E, 0x2A, 0x03, 0x04, 0x0C, 0x02,
	0x30, 0x27, 0x33, 0x14, 0x1E, 0x02, 0x04, 0x3F, 0x01, 0x1E, 0x55, 0x21,
	0x44, 0x70, 0x0B, 0x39, 0x05, 0x23, 0x12, 0x3E, 0x56, 0x25, 0x2E, 0x1B,
	0x25, 0x15, 0x14, 0x5B, 0x21, 0x3F, 0x15, 0x24, 0x20, 0x18, 0x34, 0x35,
	0x23, 0x11, 0x10, 0x58, 0x0C, 0x2D, 0x26, 0x05, 0x05, 0x58, 0x29, 0x20,
	0x06, 0x0B, 0x15, 0x17, 0x0D, 0x0C, 0x59, 0x52, 0x09, 0x2A, 0x34, 0x47,
	0x23, 0x1F, 0x3B, 0x11, 0x43, 0x58, 0x03, 0x1E, 0x03, 0x2D, 0x0A, 0x14,
	0x19, 0x04, 0x54, 0x33, 0x45, 0x5F, 0x15, 0x19, 0x02, 0x5E, 0x20, 0x0D,
	0x1F, 0x16, 0x29, 0x58, 0x0D, 0x0A, 0x22, 0x3B, 0x02, 0x73, 0x5F, 0x00,
	0x25, 0x3F, 0x04, 0x1C, 0x52, 0x2D, 0x09, 0x32, 0x2A, 0x10, 0x27, 0x05,
	0x17, 0x5B, 0x2E, 0x2B, 0x5A, 0x26, 0x1A, 0x0E, 0x0A, 0x3A, 0x06, 0x58,
	0x23, 0x0C, 0x44, 0x2F, 0x58, 0x37, 0x07, 0x59, 0x13, 0x27, 0x57, 0x00,
	0x38, 0x24, 0x5C, 0x0E, 0x19, 0x2A, 0x0F, 0x27, 0x13, 0x04, 0x5E, 0x28,
	0x19, 0x28, 0x2F, 0x5B, 0x27, 0x04, 0x54, 0x2F, 0x52, 0x0A, 0x0D, 0x0F,
	0x09, 0x3C, 0x08, 0x3C, 0x3B, 0x2F, 0x05, 0x27, 0x35, 0x32, 0x5F, 0x5B,
	0x69, 0x23, 0x09, 0x18, 0x31, 0x00, 0x22, 0x0D, 0x56, 0x19, 0x6D, 0x0B,
	0x0F, 0x38, 0x11, 0x24, 0x3D, 0x07, 0x28, 0x1B, 0x30, 0x0A, 0x19, 0x1C,
	0x3B, 0x2C, 0x2A, 0x50, 0x02, 0x1C, 0x07, 0x3D, 0x06, 0x3E, 0x40, 0x7B,
	0x16, 0x58, 0x1C, 0x33, 0x04, 0x16, 0x1B, 0x26, 0x0E, 0x04, 0x05, 0x0A,
	0x01, 0x23, 0x23, 0x28, 0x20, 0x0F, 0x33, 0x18, 0x1B, 0x36, 0x5C, 0x1D,
	0x37, 0x5B, 0x2D, 0x29, 0x2C, 0x15, 0x39, 0x30, 0x24, 0x1A, 0x75, 0x24,
	0x33, 0x22, 0x33, 0x77, 0x22, 0x16, 0x1C, 0x0E, 0x26, 0x0F, 0x0B, 0x34,
	0x06, 0x77, 0x27, 0x28, 0x18, 0x19, 0x73, 0x2A, 0x2A, 0x08, 0x29, 0x17,
	0x0A, 0x53, 0x02, 0x28, 0x23, 0x5D, 0x20, 0x3A, 0x3C, 0x2A, 0x43, 0x59,
	0x04, 0x33, 0x05, 0x1E, 0x35, 0x19, 0x31, 0x0B, 0x00, 0x54, 0x06, 0x3A,
	0x25, 0x5B, 0x2E, 0x08, 0x32, 0x75, 0x02, 0x28, 0x1C, 0x58, 0x72, 0x29,
	0x2E, 0x1E, 0x24, 0x24, 0x20, 0x29, 0x04, 0x23, 0x70, 0x38, 0x27, 0x39,
	0x13, 0x17, 0x47, 0x33, 0x56, 0x5D, 0x06, 0x00, 0x56, 0x02, 0x58, 0x72,
	0x3C, 0x29, 0x26, 0x2F, 0x34, 0x23, 0x2D, 0x59, 0x23, 0x12, 0x3D, 0x27,
	0x1C, 0x58, 0x08, 0x25, 0x33, 0x59, 0x58, 0x74, 0x05, 0x0F, 0x56, 0x39,
	0x69, 0x0E, 0x59, 0x5B, 0x39, 0x73, 0x58, 0x54, 0x5F, 0x1A, 0x00, 0x58,
	0x29, 0x45, 0x18, 0x2B, 0x5F, 0x19, 0x07, 0x04, 0x30, 0x59, 0x16, 0x28,
	0x1C, 0x21, 0x24, 0x50, 0x59, 0x05, 0x77, 0x2D, 0x27, 0x2C, 0x39, 0x71,
	0x34, 0x57, 0x3F, 0x24, 0x34, 0x5D, 0x27, 0x05, 0x32, 0x0B, 0x58, 0x2A,
	0x34, 0x0C, 0x33, 0x26, 0x2C, 0x34, 0x26, 0x27, 0x1B, 0x17, 0x25, 0x58,
	0x32, 0x03, 0x06, 0x38, 0x29, 0x7A, 0x35, 0x23, 0x19, 0x5D, 0x34, 0x1D,
	0x2F, 0x1C, 0x13, 0x2B, 0x2B, 0x12, 0x2B, 0x22, 0x2A, 0x16, 0x00, 0x56,
	0x03, 0x0D, 0x28, 0x30, 0x5C, 0x2A, 0x37, 0x38, 0x08, 0x2B, 0x3B, 0x06,
	0x34, 0x04, 0x02, 0x5B, 0x10, 0x09, 0x2C, 0x56, 0x24, 0x06, 0x03, 0x11,
	0x2D, 0x09, 0x30, 0x0D, 0x57, 0x1E, 0x28, 0x2F, 0x01, 0x08, 0x1B, 0x06,
	0x06, 0x06, 0x34, 0x01, 0x23, 0x26, 0x2D, 0x58, 0x3B, 0x3F, 0x30, 0x05,
	0x12, 0x26, 0x3A, 0x37, 0x1A, 0x37, 0x38, 0x52, 0x3A, 0x3E, 0x32, 0x23,
	0x27, 0x3B, 0x34, 0x06, 0x14, 0x1E, 0x10, 0x5E, 0x0C, 0x23, 0x28, 0x2E,
	0x26, 0x11, 0x19, 0x13, 0x29, 0x2B, 0x26, 0x14, 0x04, 0x11, 0x08, 0x0F,
	0x0D, 0x02, 0x35, 0x08, 0x17, 0x21, 0x18, 0x3A, 0x15, 0x08, 0x0F, 0x03,
	0x09, 0x19, 0x12, 0x08, 0x1C, 0x17, 0x29, 0x34, 0x08, 0x21, 0x2E, 0x36,
	0x13, 0x5E, 0x5D, 0x0E, 0x5C, 0x04, 0x24, 0x52, 0x01, 0x08, 0x54, 0x5A,
	0x38, 0x38, 0x1A, 0x4A, 0x24, 0x22, 0x33, 0x3B, 0x06, 0x5A, 0x3E, 0x7A,
	0x19, 0x07, 0x16, 0x0D, 0x04, 0x2F, 0x16, 0x59, 0x40, 0x20, 0x3B, 0x38,
	0x2A, 0x3A, 0x0E, 0x59, 0x37, 0x3A, 0x13, 0x0D, 0x35, 0x16, 0x22, 0x38,
	0x36, 0x03, 0x0C, 0x09, 0x3B, 0x1B, 0x20, 0x22, 0x3D, 0x00, 0x7B, 0x2D,
	0x2C, 0x0C, 0x2A, 0x69, 0x2A, 0x2E, 0x57, 0x32, 0x29, 0x26, 0x10, 0x0F,
	0x11, 0x32, 0x26, 0x07, 0x41, 0x39, 0x26, 0x5C, 0x15, 0x28, 0x1E, 0x13,
	0x06, 0x14, 0x39, 0x00, 0x2C, 0x5F, 0x2C, 0x2F, 0x13, 0x38, 0x3B, 0x25,
	0x59, 0x01, 0x0E, 0x27, 0x37, 0x03, 0x13, 0x0E, 0x38, 0x38, 0x20, 0x40,
	0x76, 0x5F, 0x10, 0x2F, 0x02, 0x70, 0x0A, 0x35, 0x0A, 0x3D, 0x33, 0x43,
	0x29, 0x3D, 0x1C, 0x0D, 0x14, 0x50, 0x23, 0x3B, 0x03, 0x05, 0x24, 0x2D,
	0x2D, 0x24, 0x0D, 0x0F, 0x57, 0x0D, 0x0D, 0x3F, 0x38, 0x22, 0x06, 0x7A,
	0x5B, 0x28, 0x19, 0x2F, 0x05, 0x20, 0x33, 0x34, 0x1C, 0x0E, 0x2E, 0x16,
	0x1E, 0x5B, 0x16, 0x1C, 0x2E, 0x5A, 0x0F, 0x72, 0x07, 0x13, 0x14, 0x3D,
	0x72, 0x18, 0x22, 0x1D, 0x05, 0x11, 0x2B, 0x0A, 0x09, 0x11, 0x77, 0x08,
	0x3B, 0x08, 0x24, 0x3B, 0x5E, 0x0E, 0x3A, 0x5B, 0x05, 0x18, 0x27, 0x3D,
	0x1C, 0x23, 0x54, 0x25, 0x0A, 0x3F, 0x69, 0x2D, 0x36, 0x5C, 0x09, 0x2F,
	0x24, 0x2E, 0x02, 0x19, 0x2C, 0x2B, 0x28, 0x18, 0x04, 0x06, 0x09, 0x12,
	0x5A, 0x09, 0x3A, 0x5B, 0x38, 0x2C, 0x0E, 0x69, 0x0D, 0x27, 0x38, 0x20,
	0x77, 0x19, 0x31, 0x05, 0x11, 0x29, 0x54, 0x50, 0x5A, 0x5A, 0x3A, 0x23,
	0x28, 0x08, 0x58, 0x72, 0x5B, 0x57, 0x3C, 0x09, 0x2D, 0x1E, 0x53, 0x0A,
	0x1B, 0x71, 0x19, 0x56, 0x27, 0x3F, 0x2B, 0x3C, 0x03, 0x0A, 0x40, 0x0A,
	0x1C, 0x10, 0x20, 0x5B, 0x0C, 0x29, 0x52, 0x39, 0x5F, 0x0C, 0x0B, 0x25,
	0x00, 0x1B, 0x08, 0x2F, 0x37, 0x37, 0x0E, 0x2D, 0x01, 0x11, 0x3E, 0x0E,
	0x2D, 0x01, 0x26, 0x1C, 0x0F, 0x05, 0x1A, 0x2F, 0x24, 0x0D, 0x75, 0x59,
	0x26, 0x29, 0x38, 0x01, 0x2A, 0x07, 0x0F, 0x03, 0x00, 0x02, 0x54, 0x09,
	0x2D, 0x18, 0x55, 0x0E, 0x20, 0x1C, 0x01, 0x1E, 0x39, 0x3D, 0x01, 0x3B,
	0x04, 0x32, 0x2C, 0x32, 0x70, 0x1F, 0x51, 0x5B, 0x5D, 0x0F, 0x3E, 0x55,
	0x02, 0x01, 0x09, 0x2E, 0x56, 0x3E, 0x12, 0x69, 0x24, 0x15, 0x17, 0x0C,
	0x7B, 0x5E, 0x20, 0x3F, 0x13, 0x1B, 0x0A, 0x14, 0x1D, 0x0D, 0x70, 0x08,
	0x55, 0x36, 0x3A, 0x01, 0x0D, 0x54, 0x25, 0x3E, 0x2A, 0x35, 0x24, 0x34,
	0x38, 0x2C, 0x2B, 0x56, 0x27, 0x0C, 0x69, 0x3B, 0x09, 0x2C, 0x5F, 0x10,
	0x5D, 0x02, 0x22, 0x1C, 0x7A, 0x39, 0x3B, 0x26, 0x01, 0x71, 0x3D, 0x38,
	0x04, 0x1A, 0x38, 0x08, 0x2A, 0x5F, 0x40, 0x00, 0x47, 0x03, 0x0C, 0x1E,
	0x23, 0x05, 0x39, 0x24, 0x29, 0x1A, 0x3F, 0x52, 0x5C, 0x31, 0x3B, 0x14,
	0x16, 0x3F, 0x2D, 0x7A, 0x21, 0x56, 0x5D, 0x24, 0x25, 0x3D, 0x57, 0x1E,
	0x1C, 0x0F, 0x01, 0x0A, 0x56, 0x53, 0x32, 0x29, 0x30, 0x23, 0x20, 0x2B,
	0x02, 0x2A, 0x28, 0x2C, 0x2A, 0x14, 0x05, 0x29, 0x20, 0x30, 0x3B, 0x13,
	0x45, 0x39, 0x71, 0x1F, 0x39, 0x2D, 0x27, 0x25, 0x3D, 0x34, 0x57, 0x01,
	0x36, 0x0E, 0x25, 0x16, 0x01, 0x0C, 0x0E, 0x29, 0x21, 0x00, 0x16, 0x24,
	0x58, 0x5B, 0x5C, 0x77, 0x3D, 0x0C, 0x20, 0x00, 0x2E, 0x1B, 0x33, 0x18,
	0x1F, 0x2A, 0x00, 0x57, 0x17, 0x1B, 0x21, 0x29, 0x53, 0x02, 0x2C, 0x23,
	0x2D, 0x19, 0x3D, 0x5E, 0x72, 0x1D, 0x54, 0x5B, 0x2E, 0x23, 0x19, 0x28,
	0x03, 0x59, 0x29, 0x5A, 0x31, 0x07, 0x21, 0x69, 0x01, 0x11, 0x36, 0x01,
	0x06, 0x5F, 0x30, 0x28, 0x28, 0x0F, 0x02, 0x2C, 0x07, 0x23, 0x36, 0x1C,
	0x06, 0x24, 0x2A, 0x74, 0x04, 0x17, 0x29, 0x0E, 0x38, 0x55, 0x11, 0x3C,
	0x02, 0x05, 0x04, 0x32, 0x24, 0x40, 0x09, 0x1A, 0x50, 0x5C, 0x3A, 0x06,
	0x58, 0x05, 0x01, 0x09, 0x2B, 0x5C, 0x26, 0x56, 0x2C, 0x7B, 0x24, 0x33,
	0x17, 0x09, 0x16, 0x03, 0x2D, 0x07, 0x26, 0x09, 0x14, 0x2B, 0x22, 0x1B,
	0x0F, 0x0E, 0x0B, 0x5A, 0x28, 0x01, 0x3F, 0x58, 0x41, 0x3C, 0x2A, 0x3E,
	0x0A, 0x41, 0x32, 0x2B, 0x0F, 0x4E, 0x2B, 0x1E, 0x28, 0x27, 0x39, 0x58,
	0x13, 0x26, 0x3A, 0x07, 0x27, 0x12, 0x12, 0x3A, 0x53, 0x27, 0x5F, 0x28,
	0x0A, 0x34, 0x58, 0x20, 0x3B, 0x2E, 0x50, 0x5D, 0x08, 0x0A, 0x21, 0x24,
	0x18, 0x39, 0x24, 0x27, 0x06, 0x27, 0x08, 0x00, 0x3C, 0x18, 0x5D, 0x1F,
	0x30, 0x2D, 0x4E, 0x2C, 0x1F, 0x2E, 0x5F, 0x0D, 0x0B, 0x0C, 0x69, 0x04,
	0x2F, 0x1E, 0x1F, 0x72, 0x2D, 0x20, 0x45, 0x08, 0x15, 0x2F, 0x56, 0x16,
	0x5C, 0x2A, 0x1F, 0x2B, 0x00, 0x12, 0x76, 0x1D, 0x0C, 0x16, 0x5E, 0x29,
	0x16, 0x2E, 0x02, 0x5D, 0x05, 0x1A, 0x34, 0x58, 0x03, 0x36, 0x2F, 0x20,
	0x3F, 0x53, 0x14, 0x5C, 0x1B, 0x5C, 0x05, 0x76, 0x28, 0x22, 0x25, 0x02,
	0x74, 0x2A, 0x02, 0x29, 0x24, 0x3B, 0x3E, 0x07, 0x2C, 0x22, 0x13, 0x08,
	0x0D, 0x1F, 0x20, 0x27, 0x47, 0x3B, 0x24, 0x01, 0x1B, 0x00, 0x29, 0x37,
	0x3D, 0x0E, 0x23, 0x17, 0x5A, 0x5D, 0x3B, 0x1E, 0x26, 0x16, 0x28, 0x70,
	0x21, 0x57, 0x3B, 0x5F, 0x0A, 0x55, 0x10, 0x1B, 0x25, 0x28, 0x24, 0x3B,
	0x5B, 0x2D, 0x36, 0x27, 0x2A, 0x0F, 0x22, 0x17, 0x34, 0x36, 0x38, 0x3C,
	0x34, 0x06, 0x33, 0x06, 0x0F, 0x13, 0x3B, 0x4A, 0x0D, 0x2D, 0x2B, 0x5A,
	0x4A, 0x24, 0x0F, 0x00, 0x23, 0x2F, 0x38, 0x0C, 0x23, 0x1C, 0x34, 0x0F,
	0x53, 0x1B, 0x15, 0x18, 0x5C, 0x52, 0x37, 0x27, 0x34, 0x57, 0x2A, 0x03,
	0x2F, 0x1B, 0x20, 0x26, 0x26, 0x15, 0x0D, 0x23, 0x2D, 0x34, 0x3A, 0x0C,
	0x19, 0x5A, 0x21, 0x21, 0x15, 0x5F, 0x52, 0x2F, 0x1A, 0x33, 0x28, 0x28,
	0x34, 0x0A, 0x0A, 0x5F, 0x06, 0x69, 0x05, 0x39, 0x57, 0x32, 0x2C, 0x09,
	0x09, 0x5A, 0x02, 0x0C, 0x02, 0x59, 0x0B, 0x25, 0x73, 0x19, 0x00, 0x5B,
	0x3D, 0x12, 0x2F, 0x0C, 0x1F, 0x2E, 0x69, 0x5D, 0x55, 0x14, 0x12, 0x21,
	0x16, 0x08, 0x24, 0x27, 0x70, 0x3C, 0x50, 0x36, 0x0F, 0x16, 0x59, 0x31,
	0x05, 0x5C, 0x0B, 0x24, 0x0F, 0x05, 0x5D, 0x0F, 0x58, 0x15, 0x08, 0x59,
	0x23, 0x3B, 0x2E, 0x14, 0x27, 0x7A, 0x0F, 0x56, 0x03, 0x1F, 0x2C, 0x19,
	0x14, 0x02, 0x05, 0x18, 0x54, 0x09, 0x3A, 0x12, 0x2A, 0x23, 0x0D, 0x03,
	0x5F, 0x25, 0x19, 0x37, 0x1E, 0x1F, 0x7B, 0x02, 0x12, 0x37, 0x3A, 0x20,
	0x0D, 0x0B, 0x5F, 0x5B, 0x21, 0x43, 0x2C, 0x07, 0x32, 0x25, 0x38, 0x16,
	0x3F, 0x02, 0x2E, 0x5B, 0x30, 0x29, 0x26, 0x26, 0x0B, 0x23, 0x38, 0x5F,
	0x2A, 0x21, 0x09, 0x14, 0x29, 0x06, 0x29, 0x2B, 0x18, 0x07, 0x12, 0x43,
	0x23, 0x3F, 0x3D, 0x04, 0x09, 0x34, 0x5B, 0x2A, 0x3B, 0x36, 0x0B, 0x26,
	0x5E, 0x37, 0x24, 0x15, 0x20, 0x07, 0x13, 0x3A, 0x31, 0x5E, 0x32, 0x13,
	0x03, 0x27, 0x24, 0x0C, 0x74, 0x09, 0x33, 0x0A, 0x5A, 0x73, 0x24, 0x4A,
	0x1E, 0x1F, 0x0B, 0x0F, 0x0D, 0x2B, 0x22, 0x23, 0x2E, 0x55, 0x18, 0x1B,
	0x2A, 0x16, 0x22, 0x09, 0x1A, 0x0E, 0x54, 0x50, 0x1C, 0x00, 0x26, 0x07,
	0x2F, 0x45, 0x1E, 0x06, 0x24, 0x56, 0x06, 0x1C, 0x24, 0x3F, 0x58, 0x5E,
	0x33, 0x10, 0x1E, 0x22, 0x0D, 0x58, 0x04, 0x5D, 0x2A, 0x58, 0x5C, 0x11,
	0x43, 0x23, 0x01, 0x53, 0x3A, 0x2F, 0x08, 0x1B, 0x52, 0x2A, 0x24, 0x0A,
	0x1E, 0x09, 0x2B, 0x0D, 0x29, 0x2B, 0x1D, 0x0E, 0x5C, 0x13, 0x3B, 0x59,
	0x72, 0x23, 0x2D, 0x24, 0x3A, 0x09, 0x0F, 0x15, 0x58, 0x3C, 0x11, 0x5F,
	0x17, 0x58, 0x0C, 0x21, 0x2E, 0x2D, 0x3B, 0x3F, 0x27, 0x5F, 0x10, 0x2C,
	0x28, 0x21, 0x14, 0x39, 0x22, 0x1C, 0x0F, 0x15, 0x2B, 0x19, 0x29, 0x12,
	0x2D, 0x2D, 0x2D, 0x09, 0x18, 0x00, 0x54, 0x06, 0x3A, 0x2E, 0x2E, 0x23,
	0x27, 0x1F, 0x38, 0x29, 0x39, 0x5E, 0x3D, 0x2A, 0x27, 0x59, 0x18, 0x2A,
	0x0B, 0x02, 0x39, 0x2A, 0x0C, 0x72, 0x01, 0x39, 0x2B, 0x33, 0x0D, 0x0A,
	0x35, 0x57, 0x2D, 0x38, 0x5C, 0x58, 0x39, 0x29, 0x26, 0x2F, 0x2B, 0x2B,
	0x03, 0x12, 0x24, 0x39, 0x1B, 0x02, 0x00, 0x39, 0x26, 0x03, 0x1E, 0x35,
	0x34, 0x58, 0x2F, 0x25, 0x6D, 0x01, 0x34, 0x21, 0x52, 0x69, 0x47, 0x39,
	0x5A, 0x2C, 0x18, 0x22, 0x3B, 0x3A, 0x06, 0x11, 0x0B, 0x27, 0x06, 0x31,
	0x25, 0x38, 0x4E, 0x1F, 0x13, 0x76, 0x3D, 0x19, 0x1E, 0x03, 0x2E, 0x3D,
	0x57, 0x39, 0x13, 0x32, 0x39, 0x0E, 0x3E, 0x5D, 0x15, 0x20, 0x12, 0x29,
	0x08, 0x3B, 0x34, 0x17, 0x08, 0x06, 0x72, 0x36, 0x2B, 0x00, 0x28, 0x1A,
	0x54, 0x11, 0x5A, 0x3B, 0x15, 0x54, 0x0B, 0x17, 0x20, 0x0F, 0x0A, 0x52,
	0x21, 0x5F, 0x26, 0x0E, 0x2F, 0x2B, 0x19, 0x72, 0x07, 0x18, 0x2A, 0x58,
	0x30, 0x2D, 0x18, 0x3F, 0x21, 0x3A, 0x34, 0x10, 0x2A, 0x1A, 0x75, 0x2F,
	0x2F, 0x20, 0x1B, 0x2D, 0x58, 0x35, 0x08, 0x5F, 0x00, 0x24, 0x58, 0x0C,
	0x05, 0x0E, 0x20, 0x12, 0x2B, 0x58, 0x25, 0x43, 0x2A, 0x56, 0x29, 0x7A,
	0x1B, 0x0B, 0x5F, 0x11, 0x11, 0x27, 0x2F, 0x38, 0x05, 0x15, 0x05, 0x26,
	0x16, 0x44, 0x2E, 0x03, 0x03, 0x39, 0x2E, 0x69, 0x06, 0x05, 0x41, 0x2F,
	0x21, 0x02, 0x57, 0x3B, 0x23, 0x0C, 0x25, 0x0E, 0x1C, 0x28, 0x74, 0x02,
	0x51, 0x37, 0x09, 0x1B, 0x28, 0x0E, 0x17, 0x09, 0x04, 0x06, 0x3B, 0x37,
	0x04, 0x26, 0x47, 0x23, 0x28, 0x0D, 0x0B, 0x3D, 0x08, 0x59, 0x0D, 0x0D,
	0x3E, 0x0D, 0x39, 0x32, 0x2A, 0x43, 0x2A, 0x03, 0x05, 0x72, 0x26, 0x19,
	0x01, 0x0C, 0x29, 0x08, 0x14, 0x02, 0x39, 0x06, 0x09, 0x50, 0x27, 0x52,
	0x38, 0x00, 0x2D, 0x29, 0x0F, 0x38, 0x3E, 0x2D, 0x00, 0x04, 0x24, 0x35,
	0x36, 0x1C, 0x18, 0x0D, 0x0A, 0x15, 0x0C, 0x0D, 0x0E, 0x5C, 0x09, 0x00,
	0x19, 0x0A, 0x02, 0x2C, 0x29, 0x3A, 0x3A, 0x5F, 0x4E, 0x03, 0x23, 0x35,
	0x1F, 0x10, 0x0B, 0x29, 0x12, 0x28, 0x33, 0x14, 0x2E, 0x28, 0x0D, 0x35,
	0x1B, 0x2A, 0x70, 0x08, 0x10, 0x18, 0x3F, 0x17, 0x08, 0x2A, 0x29, 0x01,
	0x07, 0x01, 0x2B, 0x2D, 0x5E, 0x11, 0x34, 0x09, 0x37, 0x5A, 0x10, 0x03,
	0x26, 0x45, 0x07, 0x76, 0x28, 0x03, 0x5C, 0x2A, 0x14, 0x3F, 0x54, 0x2C,
	0x00, 0x12, 0x59, 0x00, 0x3C, 0x5E, 0x24, 0x1A, 0x51, 0x2F, 0x53, 0x31,
	0x19, 0x57, 0x58, 0x12, 0x12, 0x03, 0x2D, 0x1C, 0x09, 0x0B, 0x19, 0x20,
	0x34, 0x44, 0x73, 0x0B, 0x2A, 0x0D, 0x5F, 0x15, 0x34, 0x2E, 0x0A, 0x01,
	0x00, 0x0F, 0x14, 0x16, 0x1B, 0x1A, 0x0A, 0x22, 0x2A, 0x28, 0x14, 0x43,
	0x09, 0x16, 0x40, 0x06, 0x5C, 0x26, 0x08, 0x5D, 0x77, 0x3F, 0x39, 0x1D,
	0x1B, 0x38, 0x01, 0x34, 0x3E, 0x5D, 0x2B, 0x43, 0x38, 0x29, 0x07, 0x26,
	0x5E, 0x12, 0x57, 0x03, 0x0D, 0x0E, 0x29, 0x23, 0x1B, 0x03, 0x16, 0x55,
	0x2B, 0x5F, 0x35, 0x3C, 0x51, 0x19, 0x07, 0x18, 0x06, 0x08, 0x5E, 0x5C,
	0x03, 0x58, 0x37, 0x26, 0x5F, 0x05, 0x0A, 0x18, 0x0F, 0x5D, 0x3A, 0x43,
	0x22, 0x0D, 0x27, 0x33, 0x24, 0x05, 0x06, 0x07, 0x35, 0x2E, 0x03, 0x1C,
	0x44, 0x07, 0x0A, 0x2A, 0x20, 0x23, 0x29, 0x5D, 0x39, 0x28, 0x04, 0x04,
	0x43, 0x13, 0x0C, 0x09, 0x11, 0x03, 0x03, 0x45, 0x0C, 0x38, 0x0D, 0x53,
	0x1C, 0x11, 0x38, 0x0F, 0x27, 0x1D, 0x11, 0x21, 0x0F, 0x20, 0x2F, 0x3D,
	0x21, 0x5E, 0x05, 0x02, 0x1B, 0x33, 0x55, 0x11, 0x2C, 0x26, 0x00, 0x38,
	0x0F, 0x02, 0x07, 0x16, 0x5D, 0x2F, 0x1E, 0x58, 0x69, 0x3B, 0x0B, 0x0D,
	0x21, 0x08, 0x3E, 0x1B, 0x21, 0x32, 0x27, 0x00, 0x0D, 0x26, 0x08, 0x2C,
	0x07, 0x2A, 0x24, 0x31, 0x35, 0x5E, 0x58, 0x23, 0x02, 0x30, 0x2A, 0x2A,
	0x21, 0x40, 0x11, 0x36, 0x23, 0x5F, 0x0A, 0x24, 0x2D, 0x26, 0x00, 0x3D,
	0x17, 0x20, 0x25, 0x08, 0x31, 0x34, 0x01, 0x00, 0x22, 0x11, 0x2F, 0x27,
	0x13, 0x2C, 0x39, 0x27, 0x2E, 0x3B, 0x41, 0x11, 0x75, 0x1A, 0x59, 0x07,
	0x13, 0x16, 0x05, 0x4E, 0x0C, 0x29, 0x2D, 0x3B, 0x0A, 0x1A, 0x08, 0x3A,
	0x19, 0x38, 0x23, 0x53, 0x2E, 0x0E, 0x2F, 0x3B, 0x53, 0x2B, 0x34, 0x4E,
	0x20, 0x2F, 0x01, 0x5B, 0x1B, 0x3B, 0x09, 0x28, 0x35, 0x27, 0x03, 0x0C,
	0x73, 0x07, 0x54, 0x0F, 0x1B, 0x11, 0x54, 0x27, 0x5C, 0x3F, 0x25, 0x25,
	0x57, 0x07, 0x1F, 0x72, 0x2A, 0x24, 0x5E, 0x0A, 0x12, 0x21, 0x55, 0x1B,
	0x05, 0x27, 0x34, 0x05, 0x29, 0x28, 0x71, 0x2F, 0x2B, 0x04, 0x53, 0x24,
	0x29, 0x2B, 0x5F, 0x5C, 0x70, 0x28, 0x0A, 0x09, 0x5E, 0x77, 0x0A, 0x53,
	0x57, 0x2F, 0x0F, 0x2F, 0x05, 0x56, 0x0C, 0x37, 0x27, 0x32, 0x25, 0x1C,
	0x0A, 0x15, 0x0B, 0x1A, 0x5F, 0x05, 0x0A, 0x56, 0x2C, 0x24, 0x77, 0x0E,
	0x54, 0x0B, 0x11, 0x38, 0x23, 0x26, 0x3E, 0x1C, 0x35, 0x21, 0x03, 0x3E,
	0x3D, 0x2F, 0x0E, 0x28, 0x3A, 0x5F, 0x75, 0x06, 0x33, 0x21, 0x08, 0x0D,
	0x0B, 0x00, 0x1B, 0x19, 0x0F, 0x20, 0x22, 0x2A, 0x44, 0x09, 0x5F, 0x34,
	0x1E, 0x2D, 0x08, 0x1C, 0x0B, 0x5C, 0x3B, 0x17, 0x55, 0x30, 0x07, 0x22,
	0x74, 0x07, 0x4E, 0x28, 0x2A, 0x2D, 0x01, 0x3B, 0x3F, 0x12, 0x11, 0x01,
	0x57, 0x37, 0x2C, 0x37, 0x24, 0x33, 0x17, 0x26, 0x0A, 0x0E, 0x50, 0x0D,
	0x5A, 0x2E, 0x1E, 0x38, 0x22, 0x02, 0x28, 0x39, 0x51, 0x59, 0x3F, 0x10,
	0x26, 0x0B, 0x56, 0x29, 0x26, 0x34, 0x57, 0x1E, 0x58, 0x2A, 0x55, 0x06,
	0x45, 0x53, 0x2D, 0x5E, 0x04, 0x3F, 0x2C, 0x70, 0x03, 0x03, 0x34, 0x1A,
	0x21, 0x39, 0x35, 0x1A, 0x2C, 0x09, 0x3C, 0x38, 0x0F, 0x1E, 0x2E, 0x54,
	0x00, 0x0F, 0x58, 0x2D, 0x5F, 0x28, 0x5F, 0x2C, 0x24, 0x23, 0x55, 0x07,
	0x38, 0x28, 0x28, 0x0E, 0x5F, 0x26, 0x0A, 0x36, 0x3B, 0x38, 0x1F, 0x01,
	0x28, 0x32, 0x01, 0x1B, 0x7A, 0x28, 0x56, 0x41, 0x26, 0x1A, 0x59, 0x0B,
	0x01, 0x0C, 0x70, 0x0B, 0x03, 0x23, 0x3C, 0x00, 0x02, 0x51, 0x2C, 0x1D,
	0x2A, 0x5D, 0x17, 0x1A, 0x07, 0x28, 0x23, 0x27, 0x20, 0x52, 0x37, 0x07,
	0x33, 0x1F, 0x01, 0x12, 0x00, 0x0F, 0x5A, 0x38, 0x1A, 0x35, 0x03, 0x1A,
	0x5B, 0x28, 0x01, 0x03, 0x3E, 0x29, 0x15, 0x35, 0x39, 0x38, 0x22, 0x0F,
	0x06, 0x0D, 0x3D, 0x21, 0x27, 0x3E, 0x57, 0x26, 0x33, 0x35, 0x58, 0x58,
	0x09, 0x38, 0x32, 0x58, 0x04, 0x3A, 0x39, 0x73, 0x5B, 0x20, 0x2C, 0x28,
	0x2B, 0x02, 0x04, 0x00, 0x22, 0x09, 0x5D, 0x2A, 0x34, 0x40, 0x07, 0x38,
	0x05, 0x3F, 0x53, 0x74, 0x01, 0x30, 0x29, 0x23, 0x69, 0x3A, 0x32, 0x20,
	0x21, 0x25, 0x25, 0x4A, 0x1C, 0x09, 0x20, 0x28, 0x24, 0x17, 0x33, 0x28,
	0x18, 0x55, 0x2A, 0x0C, 0x07, 0x09, 0x57, 0x3E, 0x59, 0x13, 0x0D, 0x26,
	0x29, 0x27, 0x29, 0x35, 0x58, 0x28, 0x19, 0x23, 0x25, 0x59, 0x09, 0x19,
	0x17, 0x16, 0x2C, 0x01, 0x2C, 0x74, 0x09, 0x32, 0x20, 0x1C, 0x12, 0x26,
	0x3B, 0x02, 0x1B, 0x31, 0x1C, 0x38, 0x5E, 0x08, 0x1B, 0x26, 0x09, 0x06,
	0x33, 0x0C, 0x04, 0x0A, 0x5E, 0x2E, 0x73, 0x36, 0x59, 0x2A, 0x11, 0x20,
	0x03, 0x25, 0x5E, 0x33, 0x09, 0x26, 0x52, 0x2B, 0x38, 0x20, 0x06, 0x1B,
	0x5D, 0x1B, 0x27, 0x2D, 0x39, 0x1A, 0x01, 0x0B, 0x1A, 0x2E, 0x2A, 0x01,
	0x06, 0x24, 0x13, 0x45, 0x0A, 0x71, 0x1B, 0x4A, 0x22, 0x3A, 0x37, 0x5A,
	0x12, 0x19, 0x1C, 0x26, 0x0E, 0x04, 0x3D, 0x53, 0x73, 0x3C, 0x24, 0x38,
	0x1F, 0x36, 0x38, 0x19, 0x2C, 0x18, 0x17, 0x1D, 0x12, 0x06, 0x5B, 0x2F,
	0x2B, 0x4A, 0x05, 0x5C, 0x01, 0x25, 0x26, 0x1E, 0x04, 0x30, 0x21, 0x2E,
	0x0C, 0x0F, 0x08, 0x1E, 0x13, 0x29, 0x03, 0x3A, 0x1D, 0x36, 0x23, 0x03,
	0x06, 0x59, 0x35, 0x2B, 0x5E, 0x3B, 0x06, 0x13, 0x05, 0x00, 0x70, 0x3D,
	0x38, 0x09, 0x3F, 0x32, 0x3D, 0x14, 0x38, 0x5B, 0x2F, 0x06, 0x15, 0x5B,
	0x09, 0x29, 0x2E, 0x57, 0x2F, 0x2C, 0x21, 0x19, 0x27, 0x5C, 0x0A, 0x37,
	0x20, 0x25, 0x3F, 0x06, 0x18, 0x03, 0x58, 0x45, 0x0D, 0x1A, 0x03, 0x06,
	0x5E, 0x27, 0x11, 0x20, 0x4A, 0x27, 0x04, 0x7A, 0x27, 0x16, 0x5D, 0x58,
	0x0F, 0x1A, 0x31, 0x0B, 0x28, 0x28, 0x2E, 0x53, 0x28, 0x1B, 0x10, 0x1A,
	0x56, 0x05, 0x1D, 0x28, 0x3F, 0x54, 0x5A, 0x26, 0x0F, 0x2E, 0x58, 0x58,
	0x52, 0x7A, 0x21, 0x23, 0x56, 0x1F, 0x32, 0x3E, 0x55, 0x03, 0x0F, 0x2B,
	0x5E, 0x2C, 0x1A, 0x2A, 0x09, 0x20, 0x57, 0x26, 0x5E, 0x2A, 0x3F, 0x07,
	0x04, 0x21, 0x69, 0x02, 0x0A, 0x14, 0x1D, 0x26, 0x25, 0x31, 0x1E, 0x0C,
	0x0B, 0x2E, 0x50, 0x1C, 0x53, 0x24, 0x29, 0x0D, 0x08, 0x09, 0x17, 0x1A,
	0x58, 0x45, 0x25, 0x32, 0x1D, 0x28, 0x58, 0x1E, 0x23, 0x43, 0x19, 0x22,
	0x1C, 0x70, 0x04, 0x17, 0x04, 0x12, 0x03, 0x08, 0x12, 0x29, 0x2C, 0x0F,
	0x3C, 0x27, 0x09, 0x31, 0x0F, 0x28, 0x55, 0x59, 0x33, 0x72, 0x20, 0x33,
	0x2D, 0x09, 0x03, 0x5A, 0x2D, 0x21, 0x40, 0x73, 0x26, 0x0F, 0x05, 0x0D,
	0x16, 0x20, 0x27, 0x16, 0x3B, 0x25, 0x1B, 0x04, 0x07, 0x2C, 0x74, 0x20,
	0x00, 0x26, 0x1F, 0x75, 0x3B, 0x54, 0x1B, 0x05, 0x23, 0x43, 0x2D, 0x27,
	0x2F, 0x08, 0x03, 0x34, 0x2B, 0x38, 0x32, 0x18, 0x03, 0x00, 0x02, 0x2D,
	0x18, 0x2E, 0x21, 0x27, 0x27, 0x58, 0x55, 0x2C, 0x06, 0x32, 0x43, 0x07,
	0x0B, 0x44, 0x38, 0x3C, 0x19, 0x3C, 0x3F, 0x6D, 0x21, 0x51, 0x3F, 0x20,
	0x18, 0x34, 0x10, 0x56, 0x06, 0x6D, 0x28, 0x0B, 0x06, 0x22, 0x08, 0x00,
	0x05, 0x41, 0x5E, 0x1B, 0x35, 0x31, 0x04, 0x5E, 0x1A, 0x16, 0x03, 0x57,
	0x03, 0x75, 0x5C, 0x31, 0x45, 0x0D, 0x29, 0x43, 0x09, 0x29, 0x1D, 0x13,
	0x1B, 0x16, 0x2B, 0x52, 0x20, 0x1E, 0x09, 0x36, 0x01, 0x05, 0x5E, 0x10,
	0x39, 0x09, 0x2B, 0x47, 0x0D, 0x5E, 0x2A, 0x1A, 0x38, 0x51, 0x5D, 0x52,
	0x0F, 0x0F, 0x04, 0x38, 0x03, 0x3B, 0x16, 0x14, 0x57, 0x09, 0x2A, 0x15,
	0x19, 0x14, 0x26, 0x25, 0x3D, 0x12, 0x19, 0x20, 0x26, 0x2D, 0x2F, 0x5D,
	0x5C, 0x6D, 0x06, 0x12, 0x1A, 0x1D, 0x73, 0x1A, 0x59, 0x08, 0x07, 0x05,
	0x09, 0x2E, 0x58, 0x0F, 0x2E, 0x35, 0x22, 0x1C, 0x3C, 0x3A, 0x54, 0x14,
	0x2A, 0x21, 0x7B, 0x1E, 0x22, 0x0D, 0x40, 0x38, 0x29, 0x2C, 0x41, 0x44,
	0x38, 0x1A, 0x23, 0x56, 0x23, 0x28, 0x5D, 0x4E, 0x03, 0x0D, 0x00, 0x54,
	0x20, 0x0B, 0x2F, 0x77, 0x21, 0x54, 0x28, 0x5F, 0x6D, 0x19, 0x25, 0x5E,
	0x5C, 0x2C, 0x04, 0x4A, 0x02, 0x5F, 0x20, 0x02, 0x17, 0x59, 0x53, 0x75,
	0x24, 0x2C, 0x41, 0x3F, 0x2C, 0x43, 0x0D, 0x06, 0x3B, 0x04, 0x43, 0x31,
	0x56, 0x23, 0x34, 0x06, 0x2F, 0x23, 0x2F, 0x34, 0x43, 0x33, 0x1E, 0x40,
	0x77, 0x15, 0x2B, 0x45, 0x5E, 0x75, 0x54, 0x2E, 0x3A, 0x52, 0x23, 0x0B,
	0x31, 0x26, 0x25, 0x24, 0x20, 0x0D, 0x45, 0x38, 0x30, 0x47, 0x31, 0x5F,
	0x26, 0x3A, 0x1C, 0x53, 0x5D, 0x0C, 0x75, 0x07, 0x13, 0x2A, 0x5D, 0x09,
	0x22, 0x19, 0x01, 0x52, 0x70, 0x2A, 0x56, 0x36, 0x3B, 0x12, 0x0F, 0x08,
	0x58, 0x28, 0x04, 0x3A, 0x4E, 0x45, 0x5E, 0x74, 0x5B, 0x03, 0x1A, 0x24,
	0x12, 0x2E, 0x02, 0x5F, 0x5F, 0x04, 0x1C, 0x57, 0x23, 0x24, 0x0A, 0x02,
	0x00, 0x02, 0x0E, 0x0B, 0x24, 0x0C, 0x1F, 0x5C, 0x0C, 0x24, 0x10, 0x01,
	0x5C, 0x2F, 0x26, 0x07, 0x02, 0x1E, 0x05, 0x34, 0x53, 0x59, 0x5D, 0x24,
	0x24, 0x10, 0x3D, 0x1D, 0x00, 0x2E, 0x22, 0x1B, 0x12, 0x01, 0x59, 0x18,
	0x2D, 0x1E, 0x37, 0x3B, 0x39, 0x5E, 0x3C, 0x08, 0x2E, 0x11, 0x37, 0x32,
	0x04, 0x28, 0x57, 0x16, 0x59, 0x2F, 0x20, 0x02, 0x3A, 0x31, 0x16, 0x27,
	0x23, 0x28, 0x0E, 0x0E, 0x09, 0x07, 0x00, 0x0C, 0x30, 0x36, 0x2E, 0x19,
	0x11, 0x05, 0x3E, 0x02, 0x0A, 0x07, 0x6D, 0x03, 0x57, 0x5F, 0x27, 0x0F,
	0x43, 0x11, 0x34, 0x04, 0x27, 0x36, 0x57, 0x34, 0x1F, 0x2C, 0x06, 0x13,
	0x1D, 0x2D, 0x21, 0x34, 0x0D, 0x0D, 0x0D, 0x35, 0x1D, 0x20, 0x22, 0x2A,
	0x26, 0x5E, 0x20, 0x37, 0x2C, 0x25, 0x0A, 0x29, 0x34, 0x52, 0x30, 0x34,
	0x11, 0x28, 0x1E, 0x24, 0x5D, 0x11, 0x2F, 0x18, 0x0F, 0x24, 0x0E, 0x57,
	0x3B, 0x00, 0x2F, 0x58, 0x16, 0x07, 0x10, 0x14, 0x0B, 0x2D, 0x5B, 0x73,
	0x3E, 0x3B, 0x16, 0x04, 0x11, 0x58, 0x50, 0x0A, 0x1E, 0x25, 0x38, 0x15,
	0x07, 0x38, 0x03, 0x2D, 0x04, 0x0A, 0x26, 0x7A, 0x16, 0x30, 0x38, 0x24,
	0x77, 0x0A, 0x2F, 0x0D, 0x07, 0x06, 0x06, 0x1B, 0x26, 0x53, 0x08, 0x3F,
	0x00, 0x21, 0x01, 0x01, 0x3D, 0x06, 0x1B, 0x3C, 0x71, 0x05, 0x37, 0x58,
	0x53, 0x72, 0x2D, 0x29, 0x06, 0x02, 0x2E, 0x22, 0x53, 0x5E, 0x39, 0x7B,
	0x54, 0x12, 0x34, 0x44, 0x01, 0x2A, 0x34, 0x5F, 0x52, 0x23, 0x34, 0x55,
	0x22, 0x1C, 0x33, 0x5F, 0x15, 0x22, 0x53, 0x13, 0x02, 0x04, 0x3D, 0x23,
	0x08, 0x34, 0x31, 0x1E, 0x39, 0x23, 0x07, 0x59, 0x5E, 0x40, 0x26, 0x1D,
	0x2F, 0x41, 0x25, 0x34, 0x47, 0x56, 0x09, 0x12, 0x3B, 0x55, 0x26, 0x36,
	0x5B, 0x05, 0x3D, 0x38, 0x5D, 0x19, 0x14, 0x1F, 0x06, 0x58, 0x1F, 0x7B,
	0x59, 0x2A, 0x1E, 0x04, 0x14, 0x14, 0x0F, 0x5D, 0x2C, 0x14, 0x0E, 0x34,
	0x28, 0x27, 0x31, 0x09, 0x2D, 0x07, 0x5A, 0x0C, 0x1D, 0x4A, 0x1E, 0x32,
	0x72, 0x20, 0x03, 0x09, 0x1C, 0x04, 0x59, 0x11, 0x34, 0x0C, 0x0F, 0x5B,
	0x02, 0x3F, 0x5A, 0x7B, 0x08, 0x13, 0x20, 0x23, 0x32, 0x39, 0x0A, 0x26,
	0x29, 0x14, 0x0A, 0x13, 0x20, 0x44, 0x35, 0x0D, 0x0D, 0x01, 0x1D, 0x2B,
	0x3D, 0x33, 0x58, 0x00, 0x28, 0x3D, 0x17, 0x2D, 0x5D, 0x2C, 0x35, 0x26,
	0x5B, 0x27, 0x2E, 0x3E, 0x3B, 0x2B, 0x07, 0x07, 0x25, 0x25, 0x1B, 0x00,
	0x20, 0x16, 0x32, 0x59, 0x00, 0x69, 0x28, 0x4E, 0x24, 0x04, 0x75, 0x36,
	0x0F, 0x1E, 0x32, 0x72, 0x25, 0x35, 0x1E, 0x3F, 0x7B, 0x05, 0x31, 0x5D,
	0x01, 0x20, 0x38, 0x2F, 0x0F, 0x5E, 0x30, 0x0F, 0x19, 0x20, 0x38, 0x35,
	0x0A, 0x23, 0x3C, 0x3C, 0x73, 0x16, 0x02, 0x17, 0x26, 0x18, 0x36, 0x52,
	0x38, 0x40, 0x01, 0x2B, 0x28, 0x58, 0x1A, 0x25, 0x22, 0x17, 0x03, 0x05,
	0x06, 0x39, 0x0E, 0x0F, 0x05, 0x36, 0x1E, 0x1B, 0x0A, 0x5B, 0x10, 0x02,
	0x50, 0x1B, 0x31, 0x76, 0x1E, 0x17, 0x2A, 0x2D, 0x04, 0x1B, 0x52, 0x23,
	0x18, 0x06, 0x24, 0x2D, 0x2D, 0x03, 0x0F, 0x1C, 0x15, 0x39, 0x09, 0x15,
	0x27, 0x0B, 0x41, 0x52, 0x0E, 0x14, 0x31, 0x0D, 0x2A, 0x38, 0x3D, 0x0C,
	0x05, 0x2C, 0x03, 0x2F, 0x54, 0x1B, 0x3E, 0x32, 0x1F, 0x23, 0x1F, 0x28,
	0x7B, 0x20, 0x0A, 0x58, 0x0C, 0x12, 0x3E, 0x29, 0x37, 0x27, 0x16, 0x15,
	0x34, 0x5D, 0x5A, 0x15, 0x35, 0x28, 0x45, 0x31, 0x73, 0x34, 0x00, 0x1E,
	0x03, 0x20, 0x02, 0x35, 0x02, 0x31, 0x3A, 0x06, 0x55, 0x59, 0x09, 0x03,
	0x26, 0x58, 0x14, 0x12, 0x2D, 0x0D, 0x23, 0x5A, 0x23, 0x04, 0x2B, 0x09,
	0x59, 0x52, 0x04, 0x3C, 0x0C, 0x16, 0x5B, 0x11, 0x43, 0x2D, 0x23, 0x53,
	0x2C, 0x0E, 0x03, 0x23, 0x28, 0x04, 0x08, 0x11, 0x5A, 0x38, 0x1B, 0x54,
	0x24, 0x1E, 0x22, 0x1A, 0x04, 0x14, 0x3F, 0x05, 0x72, 0x15, 0x27, 0x38,
	0x2E, 0x75, 0x05, 0x35, 0x5A, 0x3B, 0x37, 0x5F, 0x37, 0x39, 0x31, 0x0E,
	0x2B, 0x0B, 0x23, 0x5A, 0x10, 0x36, 0x06, 0x5A, 0x25, 0x1A, 0x0E, 0x3B,
	0x25, 0x1A, 0x31, 0x1E, 0x2C, 0x26, 0x20, 0x14, 0x5C, 0x04, 0x1F, 0x1A,
	0x18, 0x2A, 0x2C, 0x09, 0x0D, 0x21, 0x18, 0x20, 0x3A, 0x44, 0x31, 0x02,
	0x09, 0x5B, 0x3F, 0x76, 0x0F, 0x50, 0x1F, 0x02, 0x15, 0x14, 0x28, 0x1E,
	0x03, 0x69, 0x22, 0x23, 0x3F, 0x52, 0x38, 0x07, 0x12, 0x26, 0x13, 0x16,
	0x09, 0x2B, 0x2F, 0x0E, 0x33, 0x15, 0x0A, 0x2C, 0x3B, 0x1A, 0x58, 0x55,
	0x18, 0x23, 0x69, 0x2D, 0x51, 0x03, 0x07, 0x32, 0x0B, 0x50, 0x58, 0x5D,
	0x31, 0x35, 0x15, 0x57, 0x28, 0x2B, 0x5C, 0x52, 0x06, 0x1D, 0x34, 0x24,
	0x1B, 0x09, 0x05, 0x71, 0x00, 0x58, 0x36, 0x5C, 0x2E, 0x58, 0x3B, 0x03,
	0x25, 0x08, 0x38, 0x06, 0x02, 0x31, 0x2F, 0x16, 0x26, 0x0C, 0x28, 0x21,
	0x18, 0x2F, 0x01, 0x00, 0x0C, 0x15, 0x0C, 0x1D, 0x1C, 0x70, 0x04, 0x0C,
	0x00, 0x3F, 0x2A, 0x5D, 0x16, 0x0A, 0x21, 0x2B, 0x1B, 0x35, 0x1D, 0x3F,
	0x26, 0x27, 0x0C, 0x34, 0x24, 0x37, 0x03, 0x0D, 0x5D, 0x1C, 0x09, 0x0A,
	0x2F, 0x19, 0x5B, 0x0B, 0x5D, 0x10, 0x08, 0x03, 0x1A, 0x5D, 0x18, 0x1E,
	0x1C, 0x73, 0x20, 0x2F, 0x56, 0x2A, 0x7B, 0x2B, 0x08, 0x2F, 0x03, 0x2D,
	0x59, 0x32, 0x1F, 0x03, 0x71, 0x5F, 0x1B, 0x24, 0x0F, 0x13, 0x2A, 0x15,
	0x3D, 0x24, 0x32, 0x54, 0x52, 0x23, 0x1F, 0x32, 0x3A, 0x07, 0x59, 0x53,
	0x06, 0x59, 0x25, 0x05, 0x13, 0x3A, 0x29, 0x15, 0x03, 0x11, 0x06, 0x23,
	0x09, 0x58, 0x32, 0x7A, 0x0D, 0x2A, 0x1F, 0x2E, 0x17, 0x2A, 0x0D, 0x5C,
	0x2A, 0x1A, 0x19, 0x18, 0x36, 0x32, 0x7A, 0x20, 0x10, 0x39, 0x2C, 0x0B,
	0x59, 0x19, 0x04, 0x22, 0x69, 0x1F, 0x13, 0x37, 0x27, 0x69, 0x28, 0x03,
	0x22, 0x11, 0x37, 0x28, 0x26, 0x01, 0x0D, 0x69, 0x39, 0x03, 0x2D, 0x5B,
	0x69, 0x07, 0x27, 0x00, 0x29, 0x03, 0x1A, 0x30, 0x07, 0x0F, 0x7A, 0x5B,
	0x07, 0x2D, 0x2A, 0x0C, 0x0E, 0x2F, 0x05, 0x20, 0x35, 0x09, 0x14, 0x07,
	0x58, 0x21, 0x20, 0x51, 0x2D, 0x5B, 0x06, 0x0E, 0x10, 0x5F, 0x2F, 0x10,
	0x47, 0x0E, 0x3A, 0x29, 0x18, 0x38, 0x37, 0x20, 0x3D, 0x24, 0x26, 0x09,
	0x45, 0x23, 0x04, 0x00, 0x02, 0x3A, 0x0A, 0x03, 0x0B, 0x35, 0x08, 0x5E,
	0x09, 0x22, 0x16, 0x23, 0x52, 0x20, 0x07, 0x00, 0x0A, 0x0C, 0x2B, 0x19,
	0x14, 0x59, 0x0C, 0x36, 0x15, 0x2D, 0x1A, 0x1F, 0x31, 0x0B, 0x22, 0x3D,
	0x0F, 0x09, 0x5F, 0x23, 0x1B, 0x19, 0x30, 0x27, 0x0A, 0x27, 0x2E, 0x20,
	0x34, 0x28, 0x26, 0x00, 0x69, 0x34, 0x07, 0x06, 0x27, 0x2C, 0x20, 0x27,
	0x00, 0x13, 0x0A, 0x3C, 0x59, 0x19, 0x1F, 0x00, 0x1C, 0x39, 0x00, 0x59,
	0x0D, 0x3C, 0x25, 0x23, 0x20, 0x00, 0x1A, 0x14, 0x3D, 0x5B, 0x3B, 0x09,
	0x20, 0x18, 0x1B, 0x2C, 0x58, 0x22, 0x1A, 0x04, 0x7B, 0x2D, 0x2D, 0x04,
	0x21, 0x33, 0x2E, 0x32, 0x22, 0x2E, 0x69, 0x2B, 0x2C, 0x01, 0x52, 0x28,
	0x01, 0x36, 0x3E, 0x3F, 0x03, 0x2D, 0x1B, 0x2C, 0x07, 0x3B, 0x28, 0x52,
	0x2D, 0x1F, 0x09, 0x43, 0x18, 0x5C, 0x1A, 0x21, 0x2B, 0x2C, 0x14, 0x13,
	0x04, 0x3B, 0x19, 0x23, 0x3C, 0x06, 0x5C, 0x15, 0x07, 0x58, 0x74, 0x00,
	0x52, 0x5F, 0x2A, 0x08, 0x05, 0x39, 0x3B, 0x0F, 0x1A, 0x04, 0x03, 0x06,
	0x58, 0x20, 0x3D, 0x37, 0x19, 0x27, 0x25, 0x5D, 0x24, 0x1A, 0x33, 0x1A,
	0x16, 0x58, 0x38, 0x09, 0x31, 0x3F, 0x30, 0x5F, 0x26, 0x3A, 0x2F, 0x00,
	0x0F, 0x3F, 0x31, 0x2B, 0x1B, 0x0C, 0x12, 0x03, 0x16, 0x32, 0x3A, 0x44,
	0x77, 0x5C, 0x56, 0x23, 0x1D, 0x0A, 0x01, 0x0D, 0x37, 0x25, 0x0B, 0x3B,
	0x4A, 0x02, 0x1A, 0x0D, 0x0E, 0x59, 0x28, 0x58, 0x1A, 0x18, 0x22, 0x2A,
	0x25, 0x69, 0x21, 0x25, 0x16, 0x3F, 0x69, 0x55, 0x32, 0x41, 0x3B, 0x73,
	0x15, 0x31, 0x45, 0x22, 0x05, 0x1D, 0x38, 0x5C, 0x1E, 0x36, 0x0A, 0x31,
	0x45, 0x00, 0x32, 0x25, 0x27, 0x38, 0x19, 0x6D, 0x29, 0x2D, 0x59, 0x44,
	0x0D, 0x02, 0x12, 0x1A, 0x0D, 0x07, 0x09, 0x00, 0x19, 0x40, 0x00, 0x5B,
	0x20, 0x5E, 0x5A, 0x03, 0x54, 0x0E, 0x1A, 0x20, 0x05, 0x24, 0x19, 0x08,
	0x3E, 0x2C, 0x58, 0x24, 0x08, 0x2F, 0x37, 0x15, 0x14, 0x1D, 0x2E, 0x71,
	0x24, 0x0B, 0x18, 0x40, 0x6D, 0x00, 0x32, 0x2D, 0x5C, 0x6D, 0x29, 0x56,
	0x0B, 0x04, 0x1B, 0x1A, 0x09, 0x5C, 0x3E, 0x09, 0x1C, 0x4E, 0x5B, 0x0D,
	0x35, 0x18, 0x05, 0x1D, 0x44, 0x32, 0x24, 0x16, 0x41, 0x38, 0x70, 0x03,
	0x28, 0x0D, 0x04, 0x13, 0x0E, 0x22, 0x0C, 0x5E, 0x6D, 0x06, 0x15, 0x5E,
	0x40, 0x0C, 0x20, 0x39, 0x0D, 0x1D, 0x3B, 0x0E, 0x4A, 0x29, 0x5F, 0x0F,
	0x27, 0x2D, 0x58, 0x09, 0x7A, 0x35, 0x29, 0x17, 0x1E, 0x06, 0x5C, 0x32,
	0x18, 0x1A, 0x3B, 0x22, 0x29, 0x5A, 0x29, 0x34, 0x08, 0x4E, 0x1A, 0x44,
	0x08, 0x1D, 0x18, 0x01, 0x32, 0x35, 0x0F, 0x02, 0x01, 0x59, 0x0C, 0x03,
	0x2A, 0x08, 0x3A, 0x38, 0x47, 0x15, 0x24, 0x39, 0x26, 0x2B, 0x34, 0x27,
	0x32, 0x0D, 0x18, 0x18, 0x08, 0x3B, 0x04, 0x3E, 0x36, 0x1D, 0x28, 0x7A,
	0x1C, 0x15, 0x45, 0x08, 0x13, 0x09, 0x00, 0x1E, 0x05, 0x0F, 0x18, 0x27,
	0x25, 0x21, 0x29, 0x19, 0x0F, 0x58, 0x2E, 0x27, 0x1A, 0x30, 0x24, 0x1D,
	0x3A, 0x5A, 0x33, 0x27, 0x03, 0x77, 0x39, 0x25, 0x45, 0x2D, 0x2B, 0x23,
	0x4E, 0x14, 0x33, 0x70, 0x1F, 0x2B, 0x1F, 0x20, 0x06, 0x3C, 0x4E, 0x5C,
	0x25, 0x0A, 0x16, 0x16, 0x29, 0x40, 0x1B, 0x2B, 0x4E, 0x5C, 0x06, 0x0C,
	0x05, 0x1B, 0x20, 0x5F, 0x23, 0x0B, 0x17, 0x26, 0x0E, 0x09, 0x0F, 0x0F,
	0x2D, 0x25, 0x75, 0x2E, 0x2E, 0x0A, 0x22, 0x08, 0x35, 0x22, 0x1C, 0x39,
	0x0D, 0x36, 0x2D, 0x1F, 0x1C, 0x12, 0x05, 0x52, 0x05, 0x00, 0x32, 0x24,
	0x22, 0x3D, 0x1B, 0x11, 0x00, 0x23, 0x22, 0x5F, 0x26, 0x23, 0x2B, 0x39,
	0x44, 0x05, 0x0E, 0x0D, 0x2F, 0x08, 0x04, 0x5B, 0x4A, 0x5C, 0x25, 0x2C,
	0x1D, 0x3B, 0x3B, 0x5E, 0x17, 0x27, 0x15, 0x5D, 0x18, 0x12, 0x26, 0x1B,
	0x0B, 0x26, 0x29, 0x1D, 0x1B, 0x3E, 0x39, 0x2A, 0x36, 0x0D, 0x25, 0x26,
	0x00, 0x29, 0x37, 0x1E, 0x38, 0x16, 0x24, 0x09, 0x07, 0x09, 0x10, 0x3C,
	0x0A, 0x21, 0x1B, 0x35, 0x1C, 0x53, 0x07, 0x0D, 0x01, 0x03, 0x10, 0x26,
	0x02, 0x09, 0x24, 0x10, 0x3F, 0x26, 0x0C, 0x0D, 0x18, 0x2A, 0x40, 0x6D,
	0x24, 0x11, 0x1D, 0x3C, 0x1A, 0x20, 0x55, 0x23, 0x2D, 0x2F, 0x47, 0x0A,
	0x37, 0x02, 0x27, 0x5F, 0x0A, 0x28, 0x52, 0x21, 0x5B, 0x29, 0x20, 0x03,
	0x1A, 0x26, 0x22, 0x25, 0x52, 0x24, 0x47, 0x20, 0x5D, 0x5D, 0x2B, 0x2A,
	0x07, 0x2A, 0x1E, 0x7A, 0x47, 0x05, 0x27, 0x1D, 0x15, 0x27, 0x0E, 0x25,
	0x0F, 0x29, 0x23, 0x19, 0x1F, 0x04, 0x1A, 0x54, 0x12, 0x05, 0x24, 0x3A,
	0x47, 0x20, 0x3D, 0x25, 0x2D, 0x0E, 0x55, 0x1C, 0x1B, 0x14, 0x16, 0x4A,
	0x0D, 0x25, 0x24, 0x26, 0x2D, 0x1D, 0x2D, 0x18, 0x2F, 0x50, 0x36, 0x0D,
	0x09, 0x5F, 0x06, 0x5D, 0x5C, 0x09, 0x1E, 0x25, 0x21, 0x18, 0x26, 0x1F,
	0x53, 0x2B, 0x3D, 0x73, 0x0F, 0x1B, 0x39, 0x28, 0x08, 0x3F, 0x3B, 0x41,
	0x0C, 0x04, 0x3D, 0x2A, 0x36, 0x3F, 0x73, 0x5A, 0x23, 0x2F, 0x29, 0x13,
	0x08, 0x30, 0x56, 0x29, 0x2D, 0x47, 0x51, 0x27, 0x31, 0x18, 0x23, 0x36,
	0x16, 0x59, 0x1B, 0x0B, 0x37, 0x2A, 0x5D, 0x26, 0x2D, 0x56, 0x5E, 0x23,
	0x71, 0x38, 0x29, 0x45, 0x20, 0x2A, 0x0E, 0x54, 0x2B, 0x24, 0x77, 0x1B,
	0x2D, 0x0A, 0x59, 0x09, 0x5F, 0x15, 0x3D, 0x2C, 0x6D, 0x27, 0x39, 0x01,
	0x2F, 0x11, 0x1C, 0x24, 0x1B, 0x5D, 0x2D, 0x2D, 0x0D, 0x3B, 0x29, 0x77,
	0x08, 0x0F, 0x09, 0x33, 0x3A, 0x0F, 0x57, 0x3D, 0x21, 0x7B, 0x1B, 0x10,
	0x39, 0x19, 0x75, 0x06, 0x39, 0x38, 0x52, 0x05, 0x03, 0x00, 0x00, 0x1A,
	0x32, 0x28, 0x53, 0x14, 0x23, 0x37, 0x0A, 0x31, 0x27, 0x0E, 0x73, 0x38,
	0x37, 0x1B, 0x29, 0x00, 0x38, 0x50, 0x0D, 0x27, 0x18, 0x5F, 0x39, 0x38,
	0x29, 0x7A, 0x38, 0x37, 0x1E, 0x3C, 0x10, 0x24, 0x12, 0x00, 0x12, 0x75,
	0x55, 0x2D, 0x3A, 0x04, 0x20, 0x58, 0x56, 0x2A, 0x08, 0x0F, 0x08, 0x0C,
	0x20, 0x28, 0x36, 0x0A, 0x11, 0x26, 0x28, 0x32, 0x59, 0x24, 0x25, 0x05,
	0x09, 0x02, 0x05, 0x2F, 0x08, 0x6D, 0x25, 0x2C, 0x2A, 0x19, 0x27, 0x15,
	0x2B, 0x1C, 0x1A, 0x35, 0x15, 0x00, 0x3B, 0x07, 0x72, 0x2E, 0x2C, 0x36,
	0x0F, 0x34, 0x2F, 0x2A, 0x23, 0x03, 0x10, 0x09, 0x33, 0x18, 0x2F, 0x38,
	0x39, 0x4E, 0x09, 0x11, 0x74, 0x3D, 0x2B, 0x1A, 0x1E, 0x34, 0x1A, 0x38,
	0x23, 0x53, 0x7A, 0x1C, 0x36, 0x04, 0x2F, 0x2E, 0x47, 0x20, 0x5F, 0x23,
	0x01, 0x29, 0x07, 0x45, 0x38, 0x28, 0x47, 0x52, 0x22, 0x5D, 0x35, 0x02,
	0x19, 0x22, 0x06, 0x6D, 0x24, 0x09, 0x0A, 0x0E, 0x76, 0x1B, 0x37, 0x02,
	0x11, 0x69, 0x15, 0x14, 0x37, 0x21, 0x38, 0x26, 0x0D, 0x1B, 0x5F, 0x05,
	0x1A, 0x31, 0x5D, 0x03, 0x00, 0x1E, 0x19, 0x3B, 0x1C, 0x27, 0x1F, 0x0D,
	0x58, 0x53, 0x2E, 0x0B, 0x29, 0x3B, 0x52, 0x75, 0x21, 0x2E, 0x23, 0x21,
	0x77, 0x2D, 0x30, 0x3F, 0x31, 0x31, 0x01, 0x56, 0x1A, 0x3D, 0x16, 0x2E,
	0x16, 0x59, 0x5F, 0x0D, 0x23, 0x07, 0x59, 0x22, 0x1B, 0x3E, 0x32, 0x2C,
	0x33, 0x28, 0x27, 0x35, 0x05, 0x52, 0x07, 0x0E, 0x11, 0x20, 0x02, 0x71,
	0x1B, 0x3B, 0x1F, 0x23, 0x11, 0x35, 0x25, 0x28, 0x59, 0x1B, 0x04, 0x4E,
	0x22, 0x5E, 0x0A, 0x43, 0x13, 0x27, 0x08, 0x29, 0x3F, 0x37, 0x0D, 0x2D,
	0x2D, 0x2A, 0x07, 0x36, 0x31, 0x0C, 0x58, 0x1B, 0x2F, 0x1E, 0x74, 0x54,
	0x58, 0x58, 0x3C, 0x25, 0x00, 0x30, 0x06, 0x05, 0x1B, 0x3F, 0x32, 0x38,
	0x05, 0x09, 0x15, 0x02, 0x16, 0x27, 0x32, 0x47, 0x06, 0x57, 0x5A, 0x00,
	0x35, 0x54, 0x29, 0x53, 0x06, 0x18, 0x31, 0x5D, 0x29, 0x37, 0x3B, 0x14,
	0x3E, 0x00, 0x2A, 0x0B, 0x0B, 0x5A, 0x09, 0x29, 0x3E, 0x1B, 0x56, 0x11,
	0x2B, 0x19, 0x4E, 0x1D, 0x3B, 0x33, 0x59, 0x07, 0x37, 0x08, 0x21, 0x20,
	0x09, 0x1B, 0x2F, 0x0D, 0x3E, 0x07, 0x06, 0x5F, 0x24, 0x1D, 0x34, 0x0C,
	0x38, 0x15, 0x1A, 0x33, 0x26, 0x03, 0x77, 0x01, 0x0A, 0x5D, 0x39, 0x07,
	0x36, 0x54, 0x1A, 0x13, 0x18, 0x14, 0x38, 0x01, 0x5F, 0x11, 0x47, 0x22,
	0x1F, 0x11, 0x0E, 0x3B, 0x38, 0x0A, 0x07, 0x20, 0x54, 0x2A, 0x1C, 0x2F,
	0x0F, 0x05, 0x51, 0x02, 0x05, 0x75, 0x0F, 0x33, 0x22, 0x1A, 0x72, 0x2B,
	0x10, 0x2D, 0x04, 0x30, 0x59, 0x19, 0x2F, 0x1E, 0x24, 0x35, 0x33, 0x26,
	0x59, 0x0D, 0x38, 0x59, 0x5F, 0x2A, 0x38, 0x00, 0x0C, 0x3C, 0x13, 0x74,
	0x54, 0x20, 0x03, 0x40, 0x24, 0x2D, 0x18, 0x18, 0x1D, 0x20, 0x55, 0x02,
	0x06, 0x23, 0x2B, 0x0A, 0x36, 0x0D, 0x1E, 0x2C, 0x0B, 0x53, 0x58, 0x2A,
	0x09, 0x1E, 0x12, 0x00, 0x00, 0x12, 0x43, 0x0A, 0x38, 0x06, 0x3B, 0x01,
	0x2A, 0x08, 0x5A, 0x09, 0x55, 0x0D, 0x2C, 0x01, 0x35, 0x34, 0x36, 0x2D,
	0x0F, 0x73, 0x5E, 0x22, 0x03, 0x39, 0x2E, 0x05, 0x4E, 0x3D, 0x0D, 0x74,
	0x2D, 0x37, 0x5D, 0x2A, 0x16, 0x59, 0x18, 0x17, 0x2F, 0x75, 0x55, 0x53,
	0x20, 0x33, 0x05, 0x2F, 0x11, 0x5D, 0x5C, 0x04, 0x3F, 0x2E, 0x04, 0x39,
	0x21, 0x09, 0x23, 0x5C, 0x1C, 0x00, 0x2A, 0x07, 0x5C, 0x28, 0x1A, 0x25,
	0x58, 0x19, 0x3E, 0x35, 0x01, 0x3B, 0x22, 0x23, 0x00, 0x5B, 0x13, 0x21,
	0x32, 0x1A, 0x06, 0x58, 0x07, 0x13, 0x0D, 0x2F, 0x05, 0x14, 0x1F, 0x37,
	0x5D, 0x34, 0x26, 0x3D, 0x00, 0x3E, 0x4A, 0x07, 0x27, 0x32, 0x2D, 0x27,
	0x2B, 0x06, 0x13, 0x2B, 0x05, 0x2F, 0x26, 0x10, 0x03, 0x2D, 0x1B, 0x2D,
	0x16, 0x5A, 0x50, 0x17, 0x0F, 0x03, 0x34, 0x0D, 0x0C, 0x0D, 0x0B, 0x5A,
	0x00, 0x28, 0x3E, 0x69, 0x02, 0x2F, 0x27, 0x3D, 0x03, 0x24, 0x2A, 0x26,
	0x20, 0x2C, 0x22, 0x55, 0x5C, 0x13, 0x77, 0x5D, 0x25, 0x07, 0x3E, 0x38,
	0x1D, 0x37, 0x0A, 0x05, 0x26, 0x01, 0x10, 0x06, 0x3E, 0x36, 0x5B, 0x13,
	0x5E, 0x3B, 0x11, 0x19, 0x12, 0x03, 0x5C, 0x74, 0x39, 0x29, 0x08, 0x5E,
	0x07, 0x24, 0x25, 0x16, 0x19, 0x13, 0x0E, 0x34, 0x1F, 0x05, 0x23, 0x16,
	0x00, 0x0A, 0x0C, 0x24, 0x3C, 0x09, 0x23, 0x5A, 0x1B, 0x38, 0x2E, 0x2C,
	0x40, 0x3A, 0x22, 0x27, 0x5A, 0x0D, 0x23, 0x59, 0x56, 0x18, 0x25, 0x10,
	0x0B, 0x52, 0x34, 0x38, 0x10, 0x0F, 0x25, 0x20, 0x39, 0x2A, 0x28, 0x36,
	0x41, 0x0F, 0x7A, 0x35, 0x15, 0x34, 0x06, 0x18, 0x39, 0x2C, 0x1E, 0x1D,
	0x24, 0x2F, 0x23, 0x28, 0x53, 0x08, 0x54, 0x51, 0x2D, 0x0F, 0x0A, 0x26,
	0x59, 0x09, 0x00, 0x2F, 0x1A, 0x02, 0x07, 0x58, 0x36, 0x07, 0x25, 0x22,
	0x5D, 0x3A, 0x03, 0x2C, 0x45, 0x01, 0x23, 0x16, 0x16, 0x41, 0x18, 0x17,
	0x03, 0x31, 0x14, 0x38, 0x1B, 0x0D, 0x25, 0x2D, 0x32, 0x32, 0x54, 0x2E,
	0x20, 0x2C, 0x2A, 0x15, 0x2B, 0x02, 0x1B, 0x0B, 0x5C, 0x51, 0x58, 0x2E,
	0x15, 0x39, 0x08, 0x0C, 0x3F, 0x37, 0x0B, 0x36, 0x5E, 0x03, 0x34, 0x1B,
	0x03, 0x23, 0x1C, 0x15, 0x36, 0x0F, 0x5B, 0x3D, 0x3A, 0x3C, 0x35, 0x2A,
	0x2C, 0x0F, 0x18, 0x50, 0x2F, 0x08, 0x3A, 0x34, 0x25, 0x1A, 0x0E, 0x76,
	0x08, 0x23, 0x17, 0x07, 0x08, 0x2F, 0x2A, 0x58, 0x1C, 0x17, 0x5E, 0x39,
	0x29, 0x26, 0x0A, 0x1E, 0x53, 0x24, 0x26, 0x36, 0x54, 0x29, 0x41, 0x32,
	0x36, 0x5B, 0x30, 0x18, 0x40, 0x25, 0x08, 0x18, 0x0A, 0x0A, 0x09, 0x29,
	0x58, 0x06, 0x1E, 0x00, 0x0D, 0x19, 0x23, 0x1F, 0x32, 0x0F, 0x12, 0x21,
	0x3A, 0x75, 0x5E, 0x07, 0x19, 0x05, 0x30, 0x1A, 0x55, 0x2F, 0x13, 0x04,
	0x04, 0x32, 0x02, 0x39, 0x34, 0x24, 0x12, 0x0D, 0x24, 0x23, 0x39, 0x59,
	0x34, 0x09, 0x2A, 0x2B, 0x0B, 0x02, 0x12, 0x12, 0x00, 0x05, 0x0D, 0x5C,
	0x34, 0x21, 0x31, 0x0A, 0x3C, 0x04, 0x14, 0x4A, 0x5B, 0x06, 0x32, 0x01,
	0x2F, 0x3C, 0x5C, 0x30, 0x3D, 0x0B, 0x59, 0x02, 0x07, 0x5B, 0x0B, 0x39,
	0x23, 0x0F, 0x1A, 0x2E, 0x1E, 0x31, 0x7A, 0x2E, 0x23, 0x2C, 0x59, 0x3B,
	0x21, 0x30, 0x3B, 0x0F, 0x05, 0x22, 0x25, 0x45, 0x5C, 0x0F, 0x5C, 0x56,
	0x07, 0x28, 0x71, 0x1A, 0x39, 0x26, 0x04, 0x07, 0x2A, 0x13, 0x06, 0x32,
	0x23, 0x2E, 0x50, 0x1A, 0x31, 0x74, 0x5B, 0x52, 0x2A, 0x3E, 0x3B, 0x3A,
	0x05, 0x36, 0x3D, 0x0D, 0x58, 0x37, 0x57, 0x29, 0x38, 0x5F, 0x2E, 0x26,
	0x1D, 0x01, 0x3E, 0x23, 0x0A, 0x23, 0x1A, 0x2A, 0x36, 0x3E, 0x00, 0x71,
	0x27, 0x0A, 0x38, 0x33, 0x11, 0x58, 0x14, 0x38, 0x0D, 0x71, 0x5E, 0x29,
	0x5D, 0x0D, 0x72, 0x5D, 0x32, 0x57, 0x01, 0x2F, 0x07, 0x23, 0x08, 0x5B,
	0x38, 0x0E, 0x24, 0x5E, 0x53, 0x01, 0x47, 0x4E, 0x34, 0x2E, 0x06, 0x01,
	0x05, 0x3F, 0x5C, 0x76, 0x5A, 0x29, 0x23, 0x32, 0x13, 0x1E, 0x0E, 0x0F,
	0x01, 0x6D, 0x15, 0x50, 0x26, 0x18, 0x23, 0x58, 0x23, 0x21, 0x0E, 0x2B,
	0x2A, 0x55, 0x1C, 0x53, 0x21, 0x5E, 0x05, 0x28, 0x5A, 0x35, 0x59, 0x0A,
	0x17, 0x2F, 0x37, 0x2D, 0x34, 0x37, 0x05, 0x75, 0x2A, 0x23, 0x26, 0x32,
	0x2D, 0x21, 0x0B, 0x5B, 0x3E, 0x0F, 0x43, 0x08, 0x2B, 0x53, 0x14, 0x35,
	0x51, 0x0B, 0x33, 0x0A, 0x24, 0x2F, 0x00, 0x2A, 0x73, 0x5B, 0x59, 0x1D,
	0x11, 0x13, 0x24, 0x0C, 0x5D, 0x22, 0x2B, 0x00, 0x39, 0x2F, 0x5A, 0x26,
	0x3A, 0x15, 0x0A, 0x1B, 0x20, 0x1E, 0x3B, 0x1D, 0x27, 0x05, 0x3B, 0x33,
	0x03, 0x00, 0x10, 0x01, 0x00, 0x16, 0x0A, 0x2A, 0x18, 0x16, 0x2F, 0x07,
	0x29, 0x0E, 0x15, 0x0B, 0x13, 0x0F, 0x3B, 0x06, 0x3C, 0x03, 0x70, 0x2B,
	0x54, 0x56, 0x2E, 0x07, 0x3A, 0x53, 0x03, 0x18, 0x17, 0x28, 0x0C, 0x5F,
	0x03, 0x1A, 0x2D, 0x33, 0x20, 0x21, 0x32, 0x1A, 0x0C, 0x1B, 0x04, 0x73,
	0x47, 0x06, 0x14, 0x58, 0x00, 0x0F, 0x23, 0x0A, 0x0F, 0x72, 0x14, 0x53,
	0x56, 0x3E, 0x2D, 0x59, 0x57, 0x0A, 0x27, 0x16, 0x39, 0x03, 0x2B, 0x26,
	0x20, 0x28, 0x26, 0x16, 0x2C, 0x35, 0x2A, 0x17, 0x5A, 0x2F, 0x26, 0x34,
	0x4A, 0x5B, 0x5A, 0x0A, 0x1A, 0x57, 0x5A, 0x59, 0x1B, 0x43, 0x54, 0x3B,
	0x0F, 0x07, 0x1A, 0x30, 0x59, 0x00, 0x38, 0x59, 0x24, 0x45, 0x29, 0x37,
	0x07, 0x39, 0x37, 0x33, 0x29, 0x5F, 0x59, 0x3A, 0x24, 0x72, 0x24, 0x27,
	0x14, 0x18, 0x73, 0x3B, 0x53, 0x18, 0x31, 0x13, 0x00, 0x36, 0x07, 0x53,
	0x04, 0x27, 0x34, 0x1F, 0x32, 0x05, 0x59, 0x2D, 0x03, 0x5F, 0x0E, 0x5E,
	0x08, 0x3D, 0x11, 0x14, 0x5E, 0x09, 0x36, 0x3E, 0x1B, 0x58, 0x0D, 0x45,
	0x0A, 0x3A, 0x5D, 0x00, 0x5D, 0x2F, 0x05, 0x5C, 0x37, 0x07, 0x1D, 0x14,
	0x1E, 0x55, 0x29, 0x26, 0x15, 0x1D, 0x00, 0x0A, 0x2A, 0x35, 0x2A, 0x30,
	0x2A, 0x20, 0x7A, 0x5A, 0x33, 0x21, 0x0F, 0x75, 0x35, 0x2A, 0x3A, 0x53,
	0x35, 0x2F, 0x3B, 0x0D, 0x04, 0x2A, 0x1D, 0x50, 0x2B, 0x0F, 0x7A, 0x3F,
	0x10, 0x09, 0x08, 0x28, 0x2D, 0x2E, 0x09, 0x2F, 0x03, 0x35, 0x30, 0x17,
	0x12, 0x34, 0x08, 0x0A, 0x5A, 0x1C, 0x10, 0x28, 0x50, 0x59, 0x03, 0x7A,
	0x0E, 0x52, 0x2C, 0x3A, 0x30, 0x06, 0x3B, 0x2F, 0x05, 0x2E, 0x47, 0x24,
	0x2A, 0x53, 0x6D, 0x3A, 0x27, 0x1D, 0x5A, 0x75, 0x04, 0x10, 0x2F, 0x1B,
	0x77, 0x2D, 0x0A, 0x3B, 0x53, 0x7B, 0x0F, 0x56, 0x18, 0x3B, 0x0A, 0x1C,
	0x12, 0x26, 0x11, 0x2E, 0x09, 0x27, 0x0A, 0x1D, 0x0B, 0x19, 0x57, 0x5D,
	0x3E, 0x7B, 0x1F, 0x32, 0x3C, 0x22, 0x0F, 0x5E, 0x0C, 0x0D, 0x3C, 0x73,
	0x38, 0x30, 0x0F, 0x1D, 0x70, 0x14, 0x4A, 0x5C, 0x02, 0x73, 0x5C, 0x16,
	0x3A, 0x3B, 0x72, 0x08, 0x51, 0x5B, 0x08, 0x28, 0x55, 0x16, 0x39, 0x31,
	0x2D, 0x0F, 0x09, 0x06, 0x53, 0x10, 0x3A, 0x59, 0x22, 0x33, 0x33, 0x18,
	0x08, 0x5B, 0x2F, 0x71, 0x28, 0x36, 0x16, 0x5D, 0x16, 0x1E, 0x2E, 0x08,
	0x26, 0x35, 0x35, 0x25, 0x18, 0x2D, 0x20, 0x0E, 0x38, 0x38, 0x11, 0x23,
	0x2E, 0x29, 0x3E, 0x01, 0x28, 0x0D, 0x12, 0x3C, 0x59, 0x03, 0x0E, 0x26,
	0x2D, 0x12, 0x0D, 0x35, 0x31, 0x5E, 0x53, 0x32, 0x26, 0x57, 0x16, 0x1E,
	0x35, 0x16, 0x3B, 0x08, 0x1E, 0x06, 0x02, 0x12, 0x59, 0x0D, 0x09, 0x16,
	0x37, 0x58, 0x13, 0x06, 0x06, 0x07, 0x02, 0x31, 0x25, 0x00, 0x02, 0x5E,
	0x5F, 0x69, 0x5A, 0x55, 0x19, 0x24, 0x71, 0x39, 0x08, 0x07, 0x5B, 0x6D,
	0x1C, 0x2F, 0x38, 0x25, 0x2C, 0x06, 0x30, 0x28, 0x1E, 0x38, 0x3E, 0x4E,
	0x2B, 0x24, 0x2B, 0x28, 0x35, 0x5D, 0x5B, 0x2A, 0x29, 0x2C, 0x1C, 0x58,
	0x11, 0x1E, 0x15, 0x34, 0x18, 0x03, 0x5B, 0x52, 0x19, 0x1C, 0x1A, 0x08,
	0x52, 0x16, 0x29, 0x1A, 0x08, 0x10, 0x5D, 0x52, 0x0D, 0x08, 0x17, 0x06,
	0x1D, 0x24, 0x5F, 0x0C, 0x0D, 0x3E, 0x1B, 0x28, 0x54, 0x03, 0x24, 0x16,
	0x08, 0x06, 0x00, 0x38, 0x25, 0x0F, 0x50, 0x1F, 0x21, 0x77, 0x5D, 0x18,
	0x3A, 0x20, 0x0D, 0x1C, 0x06, 0x17, 0x06, 0x2A, 0x39, 0x31, 0x2F, 0x32,
	0x34, 0x2E, 0x51, 0x08, 0x3C, 0x03, 0x21, 0x29, 0x5B, 0x31, 0x15, 0x2B,
	0x2A, 0x2F, 0x1C, 0x0E, 0x58, 0x05, 0x17, 0x19, 0x0E, 0x2E, 0x53, 0x1C,
	0x1E, 0x38, 0x5B, 0x0F, 0x5D, 0x40, 0x16, 0x5A, 0x2B, 0x01, 0x1A, 0x15,
	0x36, 0x56, 0x1A, 0x5B, 0x13, 0x07, 0x30, 0x0B, 0x29, 0x00, 0x55, 0x0A,
	0x5F, 0x07, 0x08, 0x00, 0x06, 0x04, 0x26, 0x03, 0x02, 0x53, 0x36, 0x5D,
	0x04, 0x07, 0x13, 0x29, 0x1E, 0x72, 0x2A, 0x1B, 0x2A, 0x02, 0x16, 0x3C,
	0x1B, 0x3A, 0x29, 0x11, 0x2D, 0x11, 0x04, 0x5F, 0x04, 0x5B, 0x58, 0x2B,
	0x40, 0x04, 0x08, 0x0E, 0x37, 0x39, 0x70, 0x19, 0x54, 0x25, 0x0E, 0x2A,
	0x35, 0x0C, 0x5F, 0x5D, 0x3B, 0x21, 0x25, 0x17, 0x0F, 0x18, 0x21, 0x17,
	0x03, 0x2E, 0x6D, 0x1C, 0x0F, 0x2C, 0x20, 0x25, 0x15, 0x2E, 0x1D, 0x18,
	0x13, 0x16, 0x05, 0x5B, 0x1F, 0x77, 0x05, 0x0D, 0x0F, 0x33, 0x05, 0x58,
	0x25, 0x17, 0x3B, 0x73, 0x00, 0x4A, 0x5B, 0x2F, 0x13, 0x5C, 0x19, 0x5C,
	0x06, 0x09, 0x00, 0x55, 0x5A, 0x0D, 0x32, 0x19, 0x54, 0x56, 0x0D, 0x08,
	0x5E, 0x1B, 0x03, 0x0F, 0x18, 0x3B, 0x3B, 0x5D, 0x0E, 0x08, 0x47, 0x2E,
	0x0A, 0x33, 0x2A, 0x1A, 0x09, 0x24, 0x2E, 0x74, 0x21, 0x29, 0x3C, 0x5C,
	0x0F, 0x47, 0x4A, 0x0B, 0x2A, 0x15, 0x5C, 0x1B, 0x5D, 0x59, 0x37, 0x18,
	0x15, 0x41, 0x19, 0x13, 0x0B, 0x51, 0x23, 0x2C, 0x03, 0x21, 0x36, 0x23,
	0x25, 0x26, 0x20, 0x28, 0x56, 0x58, 0x0A, 0x07, 0x0D, 0x37, 0x21, 0x38,
	0x06, 0x56, 0x22, 0x02, 0x73, 0x03, 0x25, 0x1B, 0x39, 0x18, 0x3C, 0x14,
	0x21, 0x03, 0x69, 0x3A, 0x36, 0x39, 0x1E, 0x16, 0x3A, 0x10, 0x0F, 0x06,
	0x31, 0x35, 0x11, 0x01, 0x5C, 0x03, 0x2D, 0x25, 0x0C, 0x0D, 0x00, 0x34,
	0x02, 0x3E, 0x28, 0x73, 0x2F, 0x57, 0x39, 0x00, 0x0D, 0x47, 0x51, 0x37,
	0x44, 0x33, 0x2F, 0x09, 0x1A, 0x58, 0x23, 0x1B, 0x06, 0x0D, 0x3D, 0x23,
	0x2D, 0x56, 0x1B, 0x3D, 0x0B, 0x0E, 0x04, 0x29, 0x0C, 0x20, 0x35, 0x54,
	0x07, 0x1A, 0x32, 0x02, 0x52, 0x5E, 0x0E, 0x01, 0x18, 0x0D, 0x05, 0x23,
	0x75, 0x38, 0x06, 0x17, 0x2A, 0x35, 0x2A, 0x51, 0x3A, 0x5F, 0x35, 0x16,
	0x12, 0x09, 0x3B, 0x7A, 0x3E, 0x54, 0x09, 0x12, 0x27, 0x04, 0x33, 0x19,
	0x1D, 0x21, 0x27, 0x36, 0x1B, 0x02, 0x06, 0x03, 0x35, 0x3F, 0x5C, 0x31,
	0x1C, 0x19, 0x41, 0x53, 0x37, 0x16, 0x04, 0x2C, 0x3F, 0x71, 0x3F, 0x0A,
	0x19, 0x00, 0x0E, 0x5B, 0x4E, 0x3E, 0x11, 0x17, 0x2E, 0x39, 0x16, 0x02,
	0x1A, 0x19, 0x0E, 0x25, 0x1E, 0x0A, 0x1B, 0x18, 0x0A, 0x3A, 0x29, 0x59,
	0x2A, 0x3D, 0x3B, 0x00, 0x54, 0x38, 0x00, 0x33, 0x7A, 0x58, 0x0D, 0x21,
	0x20, 0x12, 0x3B, 0x2C, 0x03, 0x0F, 0x09, 0x5B, 0x51, 0x57, 0x2F, 0x33,
	0x04, 0x2F, 0x3B, 0x5C, 0x07, 0x27, 0x2D, 0x0A, 0x3D, 0x1A, 0x1A, 0x2A,
	0x3D, 0x59, 0x2B, 0x0D, 0x58, 0x1F, 0x33, 0x2F, 0x29, 0x06, 0x1F, 0x2F,
	0x15, 0x01, 0x2D, 0x3F, 0x32, 0x0E, 0x29, 0x20, 0x39, 0x23, 0x34, 0x20,
	0x20, 0x36, 0x0A, 0x7B, 0x3F, 0x25, 0x02, 0x44, 0x07, 0x16, 0x12, 0x25,
	0x0C, 0x27, 0x5F, 0x0A, 0x1E, 0x12, 0x74, 0x0B, 0x19, 0x2D, 0x20, 0x08,
	0x5C, 0x3B, 0x04, 0x1E, 0x2C, 0x07, 0x4E, 0x23, 0x5F, 0x00, 0x23, 0x0F,
	0x19, 0x08, 0x7A, 0x5C, 0x2C, 0x45, 0x0C, 0x14, 0x25, 0x24, 0x20, 0x3B,
	0x11, 0x5C, 0x27, 0x41, 0x04, 0x76, 0x1C, 0x0E, 0x1C, 0x05, 0x08, 0x0D,
	0x20, 0x09, 0x3B, 0x31, 0x22, 0x2D, 0x3E, 0x5D, 0x7A, 0x14, 0x23, 0x45,
	0x12, 0x3B, 0x36, 0x50, 0x3E, 0x5E, 0x71, 0x03, 0x17, 0x5A, 0x20, 0x2F,
	0x1A, 0x30, 0x36, 0x32, 0x18, 0x07, 0x2B, 0x36, 0x1A, 0x07, 0x5F, 0x52,
	0x2F, 0x3A, 0x70, 0x3E, 0x4A, 0x23, 0x3F, 0x7A, 0x5D, 0x29, 0x16, 0x1A,
	0x0A, 0x38, 0x56, 0x5B, 0x32, 0x30, 0x54, 0x09, 0x2D, 0x2A, 0x29, 0x03,
	0x58, 0x20, 0x26, 0x06, 0x23, 0x2F, 0x2C, 0x44, 0x32, 0x5E, 0x55, 0x19,
	0x26, 0x0C, 0x47, 0x06, 0x28, 0x0D, 0x2B, 0x23, 0x31, 0x27, 0x2E, 0x29,
	0x24, 0x30, 0x01, 0x18, 0x72, 0x1C, 0x07, 0x17, 0x07, 0x0F, 0x20, 0x16,
	0x23, 0x2E, 0x0F, 0x0A, 0x38, 0x25, 0x5F, 0x69, 0x1B, 0x26, 0x17, 0x2C,
	0x2C, 0x01, 0x08, 0x03, 0x3D, 0x12, 0x05, 0x03, 0x17, 0x2A, 0x17, 0x3B,
	0x0F, 0x37, 0x27, 0x3A, 0x3F, 0x20, 0x0F, 0x0D, 0x27, 0x2E, 0x14, 0x08,
	0x1E, 0x01, 0x15, 0x23, 0x2A, 0x38, 0x7A, 0x3B, 0x2D, 0x1D, 0x59, 0x33,
	0x23, 0x05, 0x24, 0x28, 0x70, 0x0B, 0x50, 0x08, 0x33, 0x27, 0x0F, 0x36,
	0x5A, 0x3A, 0x07, 0x5F, 0x36, 0x26, 0x18, 0x0C, 0x18, 0x14, 0x25, 0x5A,
	0x77, 0x27, 0x10, 0x3E, 0x2C, 0x26, 0x1A, 0x33, 0x3D, 0x20, 0x71, 0x0F,
	0x0D, 0x5E, 0x04, 0x2C, 0x2B, 0x00, 0x1D, 0x22, 0x15, 0x5A, 0x33, 0x17,
	0x58, 0x34, 0x5E, 0x18, 0x05, 0x32, 0x76, 0x2E, 0x51, 0x21, 0x31, 0x20,
	0x0A, 0x11, 0x34, 0x58, 0x13, 0x15, 0x10, 0x58, 0x3E, 0x0F, 0x1E, 0x3B,
	0x36, 0x23, 0x2D, 0x00, 0x0C, 0x05, 0x22, 0x12, 0x2D, 0x03, 0x3E, 0x3B,
	0x0E, 0x19, 0x13, 0x23, 0x5F, 0x0C, 0x5E, 0x13, 0x37, 0x5A, 0x2B, 0x47,
	0x50, 0x05, 0x04, 0x16, 0x03, 0x02, 0x24, 0x5F, 0x15, 0x21, 0x18, 0x0B,
	0x3F, 0x0F, 0x5D, 0x36, 0x38, 0x13, 0x2B, 0x26, 0x0F, 0x5D, 0x05, 0x1A,
	0x5C, 0x0F, 0x08, 0x1C, 0x17, 0x38, 0x39, 0x18, 0x44, 0x2E, 0x19, 0x38,
	0x08, 0x5B, 0x71, 0x3D, 0x20, 0x2F, 0x18, 0x1A, 0x0B, 0x0F, 0x58, 0x39,
	0x33, 0x5D, 0x4E, 0x23, 0x04, 0x35, 0x1A, 0x02, 0x19, 0x1B, 0x2E, 0x03,
	0x28, 0x02, 0x29, 0x69, 0x3D, 0x25, 0x2B, 0x21, 0x06, 0x03, 0x0D, 0x0C,
	0x52, 0x18, 0x3F, 0x32, 0x19, 0x27, 0x11, 0x05, 0x29, 0x28, 0x5C, 0x72,
	0x2E, 0x19, 0x21, 0x1D, 0x2C, 0x04, 0x2A, 0x05, 0x0C, 0x70, 0x04, 0x27,
	0x3C, 0x20, 0x77, 0x47, 0x36, 0x3E, 0x28, 0x24, 0x06, 0x18, 0x27, 0x3B,
	0x17, 0x23, 0x57, 0x2D, 0x22, 0x00, 0x19, 0x2D, 0x39, 0x2F, 0x08, 0x3C,
	0x0A, 0x2F, 0x40, 0x0C, 0x2D, 0x1B, 0x26, 0x0C, 0x26, 0x15, 0x57, 0x1D,
	0x1C, 0x73, 0x14, 0x19, 0x36, 0x06, 0x2D, 0x09, 0x52, 0x20, 0x0C, 0x0F,
	0x34, 0x2D, 0x2B, 0x1F, 0x04, 0x0F, 0x25, 0x3D, 0x5C, 0x37, 0x3E, 0x07,
	0x0B, 0x39, 0x75, 0x0E, 0x53, 0x3A, 0x3F, 0x30, 0x1B, 0x37, 0x0B, 0x12,
	0x06, 0x1C, 0x38, 0x41, 0x24, 0x35, 0x2B, 0x39, 0x2F, 0x2A, 0x0A, 0x1E,
	0x13, 0x3C, 0x20, 0x2E, 0x20, 0x53, 0x29, 0x5A, 0x25, 0x28, 0x3B, 0x09,
	0x28, 0x27, 0x5A, 0x31, 0x04, 0x3D, 0x01, 0x19, 0x34, 0x2D, 0x3D, 0x09,
	0x58, 0x24, 0x1E, 0x2F, 0x37, 0x39, 0x28, 0x1C, 0x18, 0x0D, 0x03, 0x0D,
	0x0D, 0x23, 0x69, 0x24, 0x37, 0x18, 0x59, 0x7B, 0x1B, 0x04, 0x1C, 0x1D,
	0x07, 0x3A, 0x00, 0x5D, 0x53, 0x38, 0x0A, 0x0B, 0x39, 0x01, 0x2F, 0x21,
	0x36, 0x1F, 0x02, 0x24, 0x1F, 0x31, 0x29, 0x19, 0x2E, 0x58, 0x58, 0x0A,
	0x3B, 0x72, 0x5F, 0x51, 0x1F, 0x44, 0x0A, 0x3D, 0x06, 0x09, 0x24, 0x15,
	0x2E, 0x14, 0x19, 0x53, 0x36, 0x0B, 0x20, 0x57, 0x23, 0x7B, 0x04, 0x1B,
	0x2D, 0x59, 0x0E, 0x5A, 0x25, 0x01, 0x1C, 0x26, 0x1F, 0x26, 0x2D, 0x3C,
	0x20, 0x29, 0x1B, 0x38, 0x3C, 0x31, 0x0B, 0x2F, 0x1A, 0x01, 0x03, 0x24,
	0x36, 0x1E, 0x0C, 0x3B, 0x00, 0x38, 0x0D, 0x3C, 0x33, 0x18, 0x29, 0x04,
	0x31, 0x2E, 0x3C, 0x0F, 0x00, 0x18, 0x24, 0x08, 0x08, 0x3D, 0x52, 0x7A,
	0x54, 0x35, 0x29, 0x26, 0x0B, 0x09, 0x0F, 0x0F, 0x26, 0x14, 0x16, 0x52,
	0x01, 0x53, 0x21, 0x1B, 0x2E, 0x57, 0x03, 0x01, 0x28, 0x0D, 0x01, 0x3E,
	0x05, 0x15, 0x57, 0x0C, 0x40, 0x04, 0x09, 0x36, 0x3B, 0x1C, 0x34, 0x0E,
	0x25, 0x14, 0x39, 0x6D, 0x18, 0x10, 0x08, 0x19, 0x20, 0x28, 0x53, 0x23,
	0x32, 0x26, 0x05, 0x50, 0x37, 0x5C, 0x28, 0x04, 0x33, 0x5A, 0x44, 0x00,
	0x29, 0x36, 0x16, 0x03, 0x2E, 0x1E, 0x20, 0x1E, 0x08, 0x09, 0x1C, 0x4E,
	0x26, 0x03, 0x05, 0x05, 0x11, 0x37, 0x5E, 0x71, 0x28, 0x00, 0x0A, 0x59,
	0x20, 0x1E, 0x17, 0x16, 0x12, 0x76, 0x09, 0x0B, 0x0C, 0x03, 0x31, 0x43,
	0x22, 0x05, 0x32, 0x3B, 0x5A, 0x15, 0x1F, 0x39, 0x28, 0x25, 0x54, 0x01,
	0x1B, 0x3B, 0x35, 0x51, 0x5C, 0x0F, 0x27, 0x21, 0x3B, 0x29, 0x0A, 0x35,
	0x24, 0x33, 0x26, 0x0A, 0x76, 0x38, 0x4E, 0x56, 0x3E, 0x36, 0x24, 0x03,
	0x5C, 0x32, 0x0F, 0x05, 0x56, 0x25, 0x09, 0x14, 0x19, 0x50, 0x41, 0x27,
	0x0E, 0x0F, 0x14, 0x34, 0x59, 0x2A, 0x43, 0x26, 0x0D, 0x44, 0x0D, 0x5D,
	0x55, 0x59, 0x06, 0x2E, 0x59, 0x52, 0x34, 0x5D, 0x05, 0x25, 0x59, 0x3F,
	0x09, 0x05, 0x0F, 0x26, 0x1A, 0x2F, 0x12, 0x00, 0x19, 0x37, 0x39, 0x0E,
	0x28, 0x53, 0x00, 0x1F, 0x04, 0x2A, 0x20, 0x59, 0x08, 0x73, 0x0F, 0x2C,
	0x45, 0x1E, 0x24, 0x58, 0x11, 0x14, 0x5D, 0x72, 0x1B, 0x29, 0x06, 0x1E,
	0x34, 0x34, 0x38, 0x56, 0x1F, 0x6D, 0x5F, 0x0E, 0x56, 0x3E, 0x35, 0x3C,
	0x15, 0x03, 0x24, 0x0A, 0x08, 0x06, 0x25, 0x40, 0x77, 0x5B, 0x58, 0x57,
	0x31, 0x10, 0x3E, 0x13, 0x34, 0x13, 0x2B, 0x59, 0x12, 0x2C, 0x12, 0x05,
	0x0B, 0x05, 0x19, 0x1E, 0x20, 0x23, 0x2D, 0x28, 0x2C, 0x11, 0x55, 0x34,
	0x07, 0x5C, 0x2A, 0x25, 0x2F, 0x19, 0x5F, 0x17, 0x1E, 0x11, 0x58, 0x00,
	0x1B, 0x0E, 0x24, 0x16, 0x1A, 0x11, 0x07, 0x4E, 0x0B, 0x00, 0x3B, 0x5E,
	0x38, 0x28, 0x1D, 0x16, 0x1F, 0x22, 0x5D, 0x05, 0x2C, 0x16, 0x56, 0x0A,
	0x59, 0x00, 0x2E, 0x31, 0x0C, 0x3C, 0x0A, 0x1F, 0x26, 0x45, 0x12, 0x18,
	0x2D, 0x27, 0x41, 0x58, 0x73, 0x39, 0x11, 0x3E, 0x31, 0x23, 0x3A, 0x2B,
	0x29, 0x22, 0x0C, 0x3C, 0x36, 0x25, 0x1C, 0x75, 0x29, 0x29, 0x1B, 0x3F,
	0x00, 0x24, 0x55, 0x0F, 0x03, 0x2B, 0x1B, 0x11, 0x3A, 0x2A, 0x00, 0x19,
	0x00, 0x1D, 0x12, 0x70, 0x39, 0x56, 0x09, 0x32, 0x18, 0x08, 0x53, 0x5A,
	0x3A, 0x0F, 0x2F, 0x50, 0x04, 0x39, 0x25, 0x29, 0x23, 0x41, 0x22, 0x69,
	0x3E, 0x56, 0x1C, 0x39, 0x2D, 0x0B, 0x0B, 0x1B, 0x2F, 0x35, 0x15, 0x29,
	0x45, 0x2E, 0x2E, 0x5A, 0x11, 0x0A, 0x0F, 0x0C, 0x2E, 0x05, 0x2B, 0x3E,
	0x2B, 0x09, 0x12, 0x1F, 0x32, 0x38, 0x5B, 0x2D, 0x1B, 0x23, 0x01, 0x01,
	0x06, 0x5C, 0x13, 0x2D, 0x28, 0x2A, 0x58, 0x5E, 0x71, 0x04, 0x0D, 0x24,
	0x06, 0x14, 0x09, 0x28, 0x04, 0x52, 0x37, 0x55, 0x2D, 0x58, 0x3F, 0x0B,
	0x19, 0x33, 0x16, 0x2C, 0x1B, 0x54, 0x15, 0x29, 0x25, 0x71, 0x3A, 0x53,
	0x25, 0x29, 0x21, 0x55, 0x53, 0x5B, 0x44, 0x2F, 0x3B, 0x25, 0x59, 0x5B,
	0x09, 0x43, 0x23, 0x5A, 0x3D, 0x1B, 0x1A, 0x0E, 0x5B, 0x2E, 0x14, 0x02,
	0x23, 0x3D, 0x3E, 0x2E, 0x29, 0x0C, 0x56, 0x21, 0x00, 0x29, 0x35, 0x18,
	0x58, 0x05, 0x2E, 0x32, 0x01, 0x03, 0x38, 0x02, 0x0B, 0x2D, 0x3F, 0x10,
	0x5E, 0x38, 0x0A, 0x59, 0x70, 0x0B, 0x13, 0x1B, 0x26, 0x20, 0x2E, 0x1B,
	0x23, 0x33, 0x0C, 0x05, 0x12, 0x3C, 0x2D, 0x30, 0x59, 0x38, 0x19, 0x2E,
	0x08, 0x1F, 0x10, 0x56, 0x00, 0x08, 0x20, 0x0B, 0x59, 0x28, 0x0D, 0x54,
	0x57, 0x34, 0x29, 0x0D, 0x0B, 0x17, 0x25, 0x26, 0x21, 0x08, 0x2F, 0x19,
	0x00, 0x70, 0x5F, 0x26, 0x3E, 0x0A, 0x35, 0x1A, 0x26, 0x23, 0x39, 0x00,
	0x01, 0x11, 0x28, 0x00, 0x74, 0x09, 0x2D, 0x36, 0x27, 0x25, 0x35, 0x26,
	0x36, 0x09, 0x13, 0x3F, 0x2E, 0x1D, 0x13, 0x75, 0x3B, 0x15, 0x1A, 0x28,
	0x0A, 0x28, 0x07, 0x41, 0x29, 0x18, 0x5F, 0x37, 0x56, 0x1E, 0x76, 0x38,
	0x54, 0x28, 0x3A, 0x06, 0x5C, 0x58, 0x3B, 0x20, 0x0B, 0x54, 0x12, 0x0B,
	0x04, 0x6D, 0x3F, 0x27, 0x5F, 0x3D, 0x30, 0x55, 0x0E, 0x01, 0x58, 0x08,
	0x1F, 0x1B, 0x04, 0x2E, 0x30, 0x54, 0x09, 0x41, 0x2A, 0x26, 0x34, 0x03,
	0x25, 0x0E, 0x31, 0x2A, 0x2E, 0x04, 0x44, 0x25, 0x27, 0x10, 0x23, 0x39,
	0x16, 0x00, 0x26, 0x21, 0x01, 0x25, 0x07, 0x24, 0x22, 0x24, 0x72, 0x2A,
	0x10, 0x18, 0x1A, 0x32, 0x02, 0x14, 0x0D, 0x38, 0x11, 0x5B, 0x26, 0x1F,
	0x1B, 0x33, 0x28, 0x30, 0x01, 0x59, 0x3B, 0x2A, 0x24, 0x1B, 0x1A, 0x23,
	0x20, 0x0F, 0x5C, 0x0F, 0x01, 0x16, 0x34, 0x5E, 0x3D, 0x2C, 0x07, 0x31,
	0x36, 0x11, 0x2F, 0x14, 0x05, 0x0D, 0x09, 0x00, 0x03, 0x00, 0x1D, 0x39,
	0x31, 0x2A, 0x52, 0x5D, 0x2A, 0x1B, 0x36, 0x4E, 0x03, 0x25, 0x32, 0x2B,
	0x0B, 0x59, 0x3B, 0x0A, 0x5C, 0x0C, 0x3E, 0x12, 0x32, 0x38, 0x18, 0x1E,
	0x3B, 0x06, 0x3B, 0x26, 0x02, 0x0E, 0x15, 0x0D, 0x17, 0x03, 0x27, 0x73,
	0x05, 0x15, 0x5A, 0x5E, 0x31, 0x0E, 0x33, 0x06, 0x1B, 0x12, 0x2A, 0x56,
	0x58, 0x40, 0x27, 0x5C, 0x02, 0x3F, 0x01, 0x3B, 0x54, 0x1B, 0x01, 0x21,
	0x23, 0x5D, 0x0A, 0x22, 0x0D, 0x38, 0x36, 0x09, 0x36, 0x1F, 0x76, 0x18,
	0x0C, 0x2D, 0x07, 0x1B, 0x3C, 0x30, 0x3A, 0x02, 0x0D, 0x03, 0x37, 0x3A,
	0x59, 0x76, 0x26, 0x19, 0x18, 0x25, 0x15, 0x08, 0x04, 0x27, 0x1E, 0x13,
	0x5F, 0x34, 0x27, 0x13, 0x38, 0x20, 0x03, 0x07, 0x27, 0x13, 0x0D, 0x0F,
	0x5C, 0x00, 0x09, 0x04, 0x0E, 0x2A, 0x5C, 0x00, 0x3B, 0x58, 0x19, 0x1F,
	0x70, 0x5C, 0x2D, 0x3C, 0x04, 0x36, 0x5B, 0x11, 0x34, 0x29, 0x72, 0x0D,
	0x0E, 0x14, 0x5F, 0x0C, 0x3C, 0x05, 0x58, 0x2E, 0x3A, 0x58, 0x08, 0x5D,
	0x3E, 0x05, 0x0B, 0x11, 0x20, 0x5E, 0x20, 0x28, 0x0E, 0x5E, 0x21, 0x20,
	0x27, 0x31, 0x1E, 0x3E, 0x03, 0x08, 0x57, 0x07, 0x0E, 0x29, 0x2B, 0x2A,
	0x07, 0x19, 0x2D, 0x3D, 0x03, 0x57, 0x2E, 0x71, 0x05, 0x07, 0x22, 0x44,
	0x33, 0x02, 0x2F, 0x24, 0x32, 0x16, 0x2D, 0x24, 0x57, 0x3C, 0x18, 0x02,
	0x0E, 0x17, 0x2F, 0x36, 0x03, 0x3B, 0x2C, 0x31, 0x27, 0x5E, 0x53, 0x39,
	0x58, 0x11, 0x18, 0x4E, 0x0F, 0x0C, 0x26, 0x00, 0x58, 0x3F, 0x06, 0x30,
	0x1D, 0x1B, 0x38, 0x1A, 0x73, 0x3D, 0x14, 0x2F, 0x13, 0x34, 0x3C, 0x12,
	0x0F, 0x2C, 0x26, 0x1A, 0x54, 0x3B, 0x28, 0x23, 0x1F, 0x17, 0x25, 0x44,
	0x7B, 0x47, 0x26, 0x20, 0x01, 0x6D, 0x21, 0x24, 0x2D, 0x01, 0x0A, 0x36,
	0x39, 0x26, 0x40, 0x32, 0x5D, 0x29, 0x34, 0x33, 0x1A, 0x29, 0x1B, 0x2C,
	0x2C, 0x0C, 0x1E, 0x17, 0x2D, 0x33, 0x06, 0x59, 0x02, 0x08, 0x2F, 0x35,
	0x35, 0x02, 0x58, 0x3C, 0x0C, 0x38, 0x4A, 0x29, 0x20, 0x38, 0x28, 0x3B,
	0x22, 0x21, 0x1A, 0x59, 0x28, 0x57, 0x00, 0x77, 0x5B, 0x2A, 0x1C, 0x53,
	0x10, 0x2A, 0x38, 0x5E, 0x44, 0x77, 0x2E, 0x4A, 0x23, 0x3B, 0x31, 0x0E,
	0x32, 0x1D, 0x0E, 0x07, 0x18, 0x2C, 0x05, 0x3E, 0x72, 0x16, 0x2D, 0x57,
	0x13, 0x10, 0x47, 0x00, 0x14, 0x04, 0x28, 0x23, 0x00, 0x1D, 0x2D, 0x6D,
	0x25, 0x0A, 0x1C, 0x5E, 0x7A, 0x54, 0x53, 0x5A, 0x5D, 0x7B, 0x2E, 0x14,
	0x24, 0x38, 0x0B, 0x38, 0x2B, 0x39, 0x0C, 0x21, 0x55, 0x30, 0x34, 0x05,
	0x38, 0x34, 0x33, 0x45, 0x32, 0x7B, 0x1B, 0x06, 0x41, 0x24, 0x24, 0x14,
	0x27, 0x3F, 0x5D, 0x71, 0x36, 0x0D, 0x3B, 0x33, 0x7B, 0x2B, 0x0A, 0x0F,
	0x1D, 0x0C, 0x59, 0x35, 0x39, 0x5E, 0x25, 0x03, 0x2E, 0x18, 0x3B, 0x15,
	0x08, 0x4A, 0x2F, 0x27, 0x0B, 0x24, 0x11, 0x56, 0x2F, 0x2C, 0x03, 0x22,
	0x41, 0x3B, 0x03, 0x0E, 0x32, 0x1C, 0x06, 0x23, 0x0D, 0x3B, 0x24, 0x13,
	0x34, 0x3D, 0x06, 0x1F, 0x3A, 0x2D, 0x5B, 0x0D, 0x0D, 0x26, 0x07, 0x5E,
	0x26, 0x28, 0x0E, 0x10, 0x24, 0x02, 0x20, 0x5C, 0x2A, 0x09, 0x0E, 0x0C,
	0x19, 0x0C, 0x08, 0x0F, 0x58, 0x5D, 0x17, 0x47, 0x36, 0x5C, 0x39, 0x7B,
	0x21, 0x2D, 0x09, 0x29, 0x15, 0x26, 0x58, 0x01, 0x0A, 0x11, 0x16, 0x38,
	0x1E, 0x1A, 0x0E, 0x43, 0x10, 0x2B, 0x59, 0x33, 0x38, 0x36, 0x41, 0x2F,
	0x08, 0x2D, 0x0A, 0x5D, 0x00, 0x71, 0x5B, 0x34, 0x3A, 0x33, 0x77, 0x47,
	0x51, 0x56, 0x28, 0x2B, 0x26, 0x0C, 0x29, 0x12, 0x0D, 0x06, 0x16, 0x1F,
	0x5B, 0x17, 0x25, 0x08, 0x17, 0x39, 0x74, 0x0E, 0x37, 0x22, 0x5F, 0x31,
	0x08, 0x08, 0x2B, 0x44, 0x0C, 0x5F, 0x56, 0x1D, 0x2D, 0x75, 0x38, 0x57,
	0x18, 0x5F, 0x77, 0x15, 0x0D, 0x38, 0x26, 0x12, 0x38, 0x0A, 0x24, 0x29,
	0x00, 0x00, 0x0B, 0x1D, 0x3B, 0x18, 0x38, 0x0A, 0x18, 0x0F, 0x2F, 0x14,
	0x52, 0x41, 0x27, 0x38, 0x58, 0x0C, 0x1F, 0x3E, 0x01, 0x1B, 0x13, 0x14,
	0x08, 0x15, 0x27, 0x29, 0x1C, 0x13, 0x3A, 0x58, 0x13, 0x03, 0x12, 0x1A,
	0x24, 0x32, 0x3C, 0x0E, 0x06, 0x27, 0x06, 0x03, 0x0F, 0x14, 0x04, 0x11,
	0x5F, 0x11, 0x30, 0x3A, 0x18, 0x2F, 0x38, 0x0F, 0x2A, 0x34, 0x3C, 0x19,
	0x05, 0x58, 0x02, 0x25, 0x3A, 0x15, 0x29, 0x32, 0x22, 0x07, 0x77, 0x07,
	0x27, 0x5C, 0x5F, 0x09, 0x38, 0x24, 0x57, 0x5B, 0x28, 0x38, 0x14, 0x0D,
	0x2F, 0x29, 0x2D, 0x09, 0x5E, 0x02, 0x08, 0x0B, 0x0C, 0x24, 0x44, 0x16,
	0x34, 0x0D, 0x26, 0x06, 0x23, 0x34, 0x03, 0x0D, 0x18, 0x05, 0x02, 0x22,
	0x0B, 0x06, 0x36, 0x3E, 0x4A, 0x5B, 0x01, 0x7A, 0x01, 0x39, 0x34, 0x5E,
	0x04, 0x06, 0x0D, 0x5C, 0x1D, 0x08, 0x2F, 0x03, 0x5A, 0x44, 0x3B, 0x2F,
	0x25, 0x1A, 0x3E, 0x1A, 0x16, 0x55, 0x57, 0x09, 0x1B, 0x1C, 0x39, 0x25,
	0x23, 0x07, 0x59, 0x2A, 0x3A, 0x3A, 0x70, 0x38, 0x2E, 0x24, 0x33, 0x24,
	0x23, 0x2A, 0x17, 0x1D, 0x71, 0x34, 0x2A, 0x56, 0x53, 0x01, 0x07, 0x59,
	0x17, 0x1B, 0x72, 0x25, 0x52, 0x5A, 0x5B, 0x36, 0x27, 0x28, 0x3B, 0x38,
	0x73, 0x1F, 0x58, 0x19, 0x13, 0x32, 0x1F, 0x2E, 0x58, 0x05, 0x11, 0x2F,
	0x35, 0x58, 0x01, 0x37, 0x24, 0x34, 0x17, 0x0D, 0x09, 0x01, 0x0E, 0x08,
	0x3D, 0x71, 0x2F, 0x05, 0x3A, 0x3D, 0x74, 0x27, 0x19, 0x58, 0x20, 0x00,
	0x05, 0x54, 0x3A, 0x31, 0x27, 0x22, 0x14, 0x5D, 0x3F, 0x10, 0x47, 0x27,
	0x56, 0x01, 0x07, 0x34, 0x15, 0x3A, 0x44, 0x04, 0x09, 0x16, 0x5B, 0x2E,
	0x2D, 0x54, 0x17, 0x23, 0x3A, 0x77, 0x16, 0x0E, 0x22, 0x22, 0x12, 0x27,
	0x2E, 0x08, 0x3A, 0x20, 0x08, 0x11, 0x58, 0x0E, 0x15, 0x03, 0x27, 0x2A,
	0x0C, 0x71, 0x36, 0x55, 0x57, 0x40, 0x36, 0x58, 0x59, 0x20, 0x5D, 0x0A,
	0x3B, 0x06, 0x28, 0x3C, 0x06, 0x3A, 0x51, 0x29, 0x3B, 0x26, 0x02, 0x2A,
	0x02, 0x0F, 0x2C, 0x3E, 0x59, 0x56, 0x2F, 0x27, 0x2E, 0x52, 0x5F, 0x26,
	0x3B, 0x19, 0x1B, 0x1E, 0x0F, 0x21, 0x2E, 0x35, 0x1B, 0x28, 0x2D, 0x15,
	0x2B, 0x5C, 0x29, 0x27, 0x5A, 0x06, 0x3F, 0x5E, 0x75, 0x02, 0x04, 0x27,
	0x0D, 0x24, 0x20, 0x59, 0x03, 0x3F, 0x15, 0x03, 0x4E, 0x3A, 0x33, 0x20,
	0x59, 0x27, 0x45, 0x0A, 0x0F, 0x5A, 0x17, 0x1A, 0x05, 0x2D, 0x2F, 0x37,
	0x28, 0x44, 0x27, 0x05, 0x2C, 0x5B, 0x2D, 0x77, 0x22, 0x28, 0x3B, 0x29,
	0x31, 0x2A, 0x2F, 0x45, 0x05, 0x10, 0x05, 0x24, 0x38, 0x18, 0x03, 0x19,
	0x15, 0x3C, 0x28, 0x2D, 0x54, 0x31, 0x3F, 0x01, 0x12, 0x55, 0x14, 0x36,
	0x3C, 0x23, 0x1A, 0x2C, 0x0D, 0x0C, 0x13, 0x16, 0x20, 0x1C, 0x04, 0x24,
	0x1B, 0x57, 0x21, 0x11, 0x0C, 0x26, 0x25, 0x56, 0x0D, 0x36, 0x35, 0x2A,
	0x37, 0x40, 0x32, 0x35, 0x2E, 0x02, 0x09, 0x29, 0x2D, 0x14, 0x5E, 0x01,
	0x35, 0x20, 0x15, 0x1C, 0x01, 0x18, 0x38, 0x15, 0x25, 0x33, 0x15, 0x26,
	0x26, 0x57, 0x38, 0x0E, 0x02, 0x35, 0x26, 0x0A, 0x03, 0x39, 0x2C, 0x1C,
	0x5C, 0x11, 0x1B, 0x54, 0x34, 0x2D, 0x34, 0x1D, 0x59, 0x5E, 0x59, 0x71,
	0x1B, 0x2D, 0x06, 0x5F, 0x38, 0x5C, 0x0A, 0x25, 0x09, 0x04, 0x28, 0x0D,
	0x1F, 0x00, 0x10, 0x18, 0x23, 0x03, 0x1A, 0x08, 0x2B, 0x18, 0x08, 0x22,
	0x0F, 0x16, 0x0D, 0x36, 0x2E, 0x74, 0x36, 0x10, 0x20, 0x53, 0x23, 0x5A,
	0x07, 0x08, 0x06, 0x28, 0x39, 0x04, 0x1A, 0x59, 0x75, 0x1E, 0x34, 0x39,
	0x2C, 0x69, 0x3C, 0x0A, 0x29, 0x31, 0x38, 0x3A, 0x02, 0x00, 0x28, 0x14,
	0x5C, 0x37, 0x3E, 0x44, 0x2B, 0x1B, 0x0E, 0x1D, 0x29, 0x10, 0x47, 0x16,
	0x3F, 0x0C, 0x1A, 0x5D, 0x37, 0x1B, 0x06, 0x25, 0x1C, 0x52, 0x59, 0x2D,
	0x7B, 0x36, 0x08, 0x24, 0x11, 0x30, 0x00, 0x39, 0x36, 0x01, 0x2F, 0x3E,
	0x53, 0x5A, 0x22, 0x0A, 0x2E, 0x23, 0x14, 0x08, 0x01, 0x3D, 0x02, 0x1D,
	0x24, 0x21, 0x1C, 0x13, 0x1D, 0x40, 0x28, 0x0B, 0x29, 0x1B, 0x22, 0x20,
	0x01, 0x12, 0x58, 0x33, 0x76, 0x1B, 0x27, 0x03, 0x2D, 0x76, 0x0E, 0x11,
	0x0D, 0x3A, 0x06, 0x1A, 0x59, 0x22, 0x20, 0x28, 0x55, 0x27, 0x5B, 0x59,
	0x14, 0x2E, 0x55, 0x0A, 0x1A, 0x20, 0x00, 0x36, 0x03, 0x11, 0x35, 0x06,
	0x38, 0x24, 0x25, 0x6D, 0x1B, 0x35, 0x00, 0x38, 0x11, 0x14, 0x50, 0x21,
	0x1D, 0x69, 0x0B, 0x59, 0x59, 0x1E, 0x00, 0x27, 0x33, 0x0A, 0x00, 0x76,
	0x1E, 0x24, 0x22, 0x11, 0x77, 0x15, 0x54, 0x0F, 0x2E, 0x16, 0x2D, 0x34,
	0x29, 0x28, 0x37, 0x15, 0x20, 0x16, 0x06, 0x76, 0x35, 0x18, 0x0A, 0x32,
	0x23, 0x0B, 0x10, 0x0F, 0x12, 0x1A, 0x00, 0x1B, 0x21, 0x1F, 0x16, 0x02,
	0x59, 0x05, 0x08, 0x2A, 0x23, 0x27, 0x0B, 0x3B, 0x13, 0x24, 0x22, 0x39,
	0x2E, 0x17, 0x0F, 0x4A, 0x24, 0x2E, 0x32, 0x5D, 0x06, 0x29, 0x0A, 0x09,
	0x0D, 0x33, 0x0F, 0x0E, 0x12, 0x07, 0x0E, 0x2C, 0x26, 0x2D, 0x09, 0x2B,
	0x20, 0x3E, 0x3A, 0x5A, 0x0C, 0x26, 0x0D, 0x71, 0x06, 0x32, 0x25, 0x13,
	0x0A, 0x21, 0x31, 0x3A, 0x2A, 0x06, 0x2F, 0x26, 0x3C, 0x44, 0x21, 0x03,
	0x2E, 0x28, 0x0E, 0x2B, 0x3F, 0x10, 0x34, 0x0F, 0x0E, 0x22, 0x28, 0x18,
	0x0C, 0x2F, 0x05, 0x4A, 0x3F, 0x00, 0x24, 0x16, 0x28, 0x09, 0x58, 0x0C,
	0x1B, 0x58, 0x20, 0x5A, 0x31, 0x24, 0x34, 0x38, 0x33, 0x26, 0x23, 0x09,
	0x02, 0x3D, 0x28, 0x3B, 0x18, 0x1E, 0x5A, 0x31, 0x00, 0x02, 0x5E, 0x0F,
	0x23, 0x59, 0x34, 0x08, 0x5F, 0x77, 0x28, 0x4A, 0x59, 0x18, 0x2C, 0x29,
	0x38, 0x5F, 0x24, 0x01, 0x1E, 0x0C, 0x37, 0x5D, 0x77, 0x21, 0x36, 0x1E,
	0x0C, 0x12, 0x01, 0x37, 0x2A, 0x1E, 0x2F, 0x1B, 0x02, 0x1A, 0x52, 0x0F,
	0x18, 0x26, 0x5E, 0x11, 0x11, 0x1A, 0x00, 0x17, 0x38, 0x05, 0x0E, 0x36,
	0x57, 0x2E, 0x0C, 0x5E, 0x04, 0x34, 0x27, 0x04, 0x58, 0x05, 0x17, 0x2D,
	0x2B, 0x43, 0x05, 0x06, 0x3C, 0x2D, 0x2D, 0x23, 0x34, 0x0A, 0x77, 0x28,
	0x04, 0x38, 0x03, 0x27, 0x01, 0x03, 0x1E, 0x2E, 0x26, 0x23, 0x56, 0x24,
	0x5E, 0x28, 0x0F, 0x04, 0x19, 0x28, 0x73, 0x35, 0x13, 0x1A, 0x33, 0x0D,
	0x08, 0x3B, 0x2B, 0x05, 0x31, 0x38, 0x2B, 0x19, 0x21, 0x28, 0x1F, 0x35,
	0x05, 0x2A, 0x23, 0x1A, 0x51, 0x0D, 0x08, 0x17, 0x35, 0x2C, 0x16, 0x0F,
	0x17, 0x1E, 0x54, 0x2A, 0x0E, 0x21, 0x36, 0x3B, 0x22, 0x40, 0x01, 0x0D,
	0x2F, 0x39, 0x12, 0x08, 0x3D, 0x34, 0x03, 0x0F, 0x23, 0x3D, 0x08, 0x0B,
	0x05, 0x21, 0x3B, 0x53, 0x58, 0x27, 0x25, 0x0F, 0x14, 0x0C, 0x19, 0x7B,
	0x36, 0x25, 0x07, 0x29, 0x29, 0x43, 0x28, 0x45, 0x33, 0x0C, 0x24, 0x1B,
	0x3E, 0x07, 0x3A, 0x1A, 0x0E, 0x1C, 0x1C, 0x12, 0x05, 0x38, 0x3C, 0x04,
	0x73, 0x19, 0x2B, 0x01, 0x12, 0x34, 0x1B, 0x16, 0x26, 0x26, 0x0C, 0x02,
	0x37, 0x06, 0x02, 0x34, 0x2E, 0x59, 0x24, 0x1E, 0x14, 0x18, 0x24, 0x16,
	0x2A, 0x24, 0x2A, 0x12, 0x27, 0x11, 0x24, 0x1C, 0x2E, 0x0A, 0x5C, 0x7B,
	0x0D, 0x1B, 0x16, 0x21, 0x7A, 0x0B, 0x17, 0x1B, 0x31, 0x75, 0x15, 0x56,
	0x2D, 0x2F, 0x26, 0x21, 0x30, 0x56, 0x2F, 0x75, 0x3C, 0x10, 0x58, 0x03,
	0x75, 0x01, 0x0A, 0x3E, 0x19, 0x2C, 0x1F, 0x20, 0x16, 0x2A, 0x13, 0x2F,
	0x0E, 0x00, 0x1E, 0x6D, 0x2E, 0x12, 0x3F, 0x13, 0x74, 0x1F, 0x00, 0x1B,
	0x00, 0x0A, 0x54, 0x27, 0x09, 0x1B, 0x03, 0x1F, 0x39, 0x0C, 0x28, 0x07,
	0x39, 0x19, 0x3F, 0x2A, 0x75, 0x38, 0x14, 0x1E, 0x3E, 0x2A, 0x5C, 0x2F,
	0x25, 0x5E, 0x08, 0x23, 0x2E, 0x39, 0x18, 0x3A, 0x24, 0x2E, 0x09, 0x59,
	0x26, 0x0B, 0x09, 0x18, 0x24, 0x09, 0x35, 0x0D, 0x1A, 0x59, 0x74, 0x43,
	0x0B, 0x1B, 0x38, 0x0D, 0x21, 0x16, 0x25, 0x0E, 0x14, 0x2E, 0x15, 0x06,
	0x00, 0x35, 0x1C, 0x0B, 0x0C, 0x0F, 0x08, 0x16, 0x02, 0x0F, 0x29, 0x03,
	0x25, 0x51, 0x1B, 0x25, 0x07, 0x27, 0x24, 0x37, 0x23, 0x6D, 0x01, 0x2C,
	0x0D, 0x38, 0x76, 0x0B, 0x11, 0x0B, 0x2E, 0x0E, 0x15, 0x0B, 0x2C, 0x25,
	0x14, 0x0B, 0x07, 0x39, 0x33, 0x0D, 0x2E, 0x25, 0x0C, 0x52, 0x35, 0x5C,
	0x53, 0x09, 0x27, 0x24, 0x05, 0x0C, 0x0A, 0x12, 0x00, 0x34, 0x0D, 0x17,
	0x58, 0x71, 0x20, 0x02, 0x14, 0x5E, 0x2D, 0x16, 0x29, 0x23, 0x3B, 0x1A,
	0x3C, 0x2B, 0x03, 0x0A, 0x3A, 0x19, 0x2D, 0x59, 0x00, 0x7B, 0x18, 0x2A,
	0x0F, 0x11, 0x01, 0x47, 0x4E, 0x45, 0x59, 0x25, 0x1F, 0x10, 0x26, 0x21,
	0x2F, 0x5A, 0x12, 0x2B, 0x21, 0x15, 0x5F, 0x37, 0x17, 0x39, 0x38, 0x1C,
	0x0D, 0x22, 0x1A, 0x0F, 0x47, 0x25, 0x18, 0x11, 0x14, 0x59, 0x38, 0x1E,
	0x19, 0x2F, 0x5C, 0x37, 0x3A, 0x29, 0x34, 0x21, 0x26, 0x0D, 0x12, 0x21,
	0x21, 0x09, 0x00, 0x20, 0x25, 0x5A, 0x32, 0x26, 0x26, 0x7A, 0x38, 0x19,
	0x00, 0x04, 0x2C, 0x07, 0x31, 0x2F, 0x22, 0x2D, 0x54, 0x23, 0x23, 0x5D,
	0x0F, 0x5B, 0x09, 0x22, 0x06, 0x71, 0x5C, 0x03, 0x5F, 0x5F, 0x77, 0x00,
	0x09, 0x19, 0x1A, 0x76, 0x16, 0x57, 0x59, 0x21, 0x0E, 0x58, 0x1B, 0x1F,
	0x25, 0x37, 0x25, 0x19, 0x2B, 0x12, 0x13, 0x34, 0x31, 0x2F, 0x1A, 0x0D,
	0x34, 0x52, 0x1C, 0x40, 0x3B, 0x03, 0x39, 0x27, 0x22, 0x03, 0x3F, 0x38,
	0x3B, 0x0C, 0x13, 0x5C, 0x2B, 0x1A, 0x3E, 0x0C, 0x5E, 0x54, 0x45, 0x29,
	0x08, 0x35, 0x28, 0x5C, 0x24, 0x25, 0x58, 0x13, 0x2A, 0x3A, 0x27, 0x36,
	0x0A, 0x07, 0x59, 0x25, 0x5F, 0x52, 0x2B, 0x59, 0x2D, 0x03, 0x0C, 0x41,
	0x13, 0x11, 0x14, 0x08, 0x03, 0x24, 0x31, 0x23, 0x23, 0x1B, 0x3C, 0x12,
	0x1F, 0x29, 0x0C, 0x1B, 0x2C, 0x3C, 0x10, 0x36, 0x01, 0x34, 0x28, 0x54,
	0x37, 0x5B, 0x16, 0x0B, 0x0B, 0x1B, 0x21, 0x01, 0x1F, 0x56, 0x02, 0x1B,
	0x06, 0x22, 0x29, 0x28, 0x0F, 0x38, 0x1E, 0x14, 0x5C, 0x5D, 0x16, 0x5E,
	0x03, 0x06, 0x3A, 0x2A, 0x1D, 0x36, 0x01, 0x3F, 0x73, 0x20, 0x28, 0x0B,
	0x0D, 0x20, 0x03, 0x0E, 0x17, 0x20, 0x01, 0x16, 0x51, 0x07, 0x0A, 0x34,
	0x3D, 0x0B, 0x0F, 0x2D, 0x28, 0x27, 0x17, 0x2D, 0x0A, 0x0F, 0x1B, 0x30,
	0x25, 0x0D, 0x33, 0x07, 0x02, 0x38, 0x11, 0x16, 0x3D, 0x2B, 0x22, 0x3F,
	0x2C, 0x26, 0x39, 0x5E, 0x01, 0x33, 0x22, 0x52, 0x00, 0x1D, 0x33, 0x2F,
	0x59, 0x5B, 0x02, 0x77, 0x0E, 0x55, 0x03, 0x5C, 0x04, 0x1E, 0x06, 0x03,
	0x1B, 0x21, 0x1F, 0x25, 0x3B, 0x3C, 0x0F, 0x1A, 0x16, 0x3C, 0x3C, 0x20,
	0x09, 0x37, 0x20, 0x22, 0x71, 0x5A, 0x17, 0x5B, 0x0C, 0x3A, 0x38, 0x0F,
	0x29, 0x08, 0x29, 0x2A, 0x27, 0x03, 0x3D, 0x0F, 0x29, 0x25, 0x5D, 0x03,
	0x33, 0x16, 0x55, 0x2C, 0x0F, 0x70, 0x5F, 0x23, 0x5F, 0x52, 0x08, 0x09,
	0x1B, 0x0C, 0x3E, 0x27, 0x21, 0x25, 0x38, 0x23, 0x2C, 0x1D, 0x03, 0x02,
	0x04, 0x76, 0x05, 0x26, 0x0F, 0x0D, 0x16, 0x01, 0x58, 0x37, 0x2C, 0x30,
	0x1A, 0x26, 0x07, 0x2A, 0x11, 0x36, 0x51, 0x04, 0x58, 0x11, 0x09, 0x0A,
	0x38, 0x58, 0x08, 0x5D, 0x59, 0x20, 0x27, 0x14, 0x29, 0x12, 0x1B, 0x44,
	0x28, 0x22, 0x27, 0x17, 0x5F, 0x06, 0x1D, 0x1B, 0x38, 0x1F, 0x30, 0x02,
	0x2A, 0x01, 0x5A, 0x73, 0x09, 0x2E, 0x3E, 0x5F, 0x0A, 0x2F, 0x0A, 0x1B,
	0x2D, 0x37, 0x5F, 0x20, 0x58, 0x06, 0x07, 0x29, 0x57, 0x41, 0x1B, 0x0C,
	0x35, 0x4E, 0x3B, 0x13, 0x25, 0x5F, 0x08, 0x41, 0x29, 0x0F, 0x0D, 0x58,
	0x00, 0x3D, 0x2E, 0x59, 0x15, 0x0F, 0x3E, 0x04, 0x14, 0x12, 0x5D, 0x3C,
	0x11, 0x20, 0x36, 0x34, 0x0A, 0x0F, 0x2E, 0x06, 0x02, 0x1C, 0x31, 0x59,
	0x0B, 0x20, 0x1D, 0x72, 0x19, 0x27, 0x39, 0x0E, 0x03, 0x54, 0x17, 0x3A,
	0x08, 0x23, 0x38, 0x2C, 0x20, 0x5F, 0x21, 0x3F, 0x3B, 0x0F, 0x04, 0x06,
	0x5E, 0x18, 0x05, 0x2C, 0x08, 0x1B, 0x16, 0x0F, 0x11, 0x38, 0x1F, 0x09,
	0x22, 0x12, 0x17, 0x09, 0x35, 0x28, 0x28, 0x00, 0x5C, 0x30, 0x27, 0x1D,
	0x14, 0x19, 0x2A, 0x00, 0x22, 0x38, 0x08, 0x09, 0x04, 0x2D, 0x1B, 0x1E,
	0x38, 0x45, 0x3E, 0x01, 0x1F, 0x10, 0x20, 0x3B, 0x03, 0x23, 0x10, 0x2D,
	0x0C, 0x31, 0x22, 0x38, 0x03, 0x1A, 0x76, 0x18, 0x28, 0x24, 0x26, 0x33,
	0x5D, 0x11, 0x56, 0x2F, 0x34, 0x2E, 0x52, 0x17, 0x31, 0x00, 0x2B, 0x16,
	0x09, 0x23, 0x08, 0x27, 0x00, 0x2B, 0x00, 0x30, 0x3C, 0x2F, 0x0D, 0x31,
	0x06, 0x35, 0x25, 0x05, 0x00, 0x3A, 0x14, 0x32, 0x1B, 0x12, 0x2B, 0x04,
	0x38, 0x3F, 0x58, 0x2A, 0x1E, 0x04, 0x0B, 0x19, 0x72, 0x25, 0x57, 0x0D,
	0x3B, 0x70, 0x3B, 0x31, 0x17, 0x2D, 0x21, 0x2E, 0x4A, 0x2A, 0x2D, 0x08,
	0x1A, 0x03, 0x0A, 0x3D, 0x32, 0x5B, 0x4E, 0x56, 0x3B, 0x7B, 0x23, 0x00,
	0x57, 0x3A, 0x2B, 0x18, 0x37, 0x2C, 0x3E, 0x05, 0x18, 0x0C, 0x14, 0x13,
	0x2C, 0x18, 0x0D, 0x5A, 0x02, 0x32, 0x0A, 0x26, 0x3A, 0x13, 0x31, 0x5C,
	0x54, 0x2D, 0x59, 0x21, 0x3B, 0x36, 0x41, 0x0F, 0x28, 0x1E, 0x58, 0x25,
	0x52, 0x03, 0x0B, 0x36, 0x27, 0x40, 0x24, 0x1E, 0x27, 0x1C, 0x5B, 0x13,
	0x24, 0x0B, 0x3D, 0x3D, 0x7A, 0x2E, 0x2C, 0x2D, 0x00, 0x07, 0x5A, 0x30,
	0x1E, 0x58, 0x04, 0x0A, 0x3B, 0x14, 0x32, 0x74, 0x35, 0x16, 0x08, 0x32,
	0x13, 0x19, 0x08, 0x5B, 0x28, 0x28, 0x08, 0x2F, 0x08, 0x40, 0x33, 0x2A,
	0x0A, 0x22, 0x5D, 0x06, 0x23, 0x37, 0x08, 0x09, 0x11, 0x39, 0x31, 0x3F,
	0x5D, 0x18, 0x0E, 0x26, 0x58, 0x1B, 0x00, 0x24, 0x52, 0x45, 0x3B, 0x0A,
	0x5C, 0x03, 0x5A, 0x13, 0x04, 0x23, 0x0A, 0x39, 0x5B, 0x70, 0x00, 0x0B,
	0x2A, 0x0C, 0x70, 0x28, 0x32, 0x26, 0x1F, 0x7A, 0x1B, 0x07, 0x19, 0x31,
	0x0E, 0x5A, 0x27, 0x1E, 0x20, 0x75, 0x5D, 0x32, 0x5B, 0x23, 0x1B, 0x25,
	0x2E, 0x23, 0x5F, 0x21, 0x5A, 0x3B, 0x22, 0x0A, 0x34, 0x59, 0x2F, 0x5F,
	0x27, 0x10, 0x5A, 0x57, 0x3C, 0x01, 0x05, 0x2E, 0x24, 0x2B, 0x00, 0x03,
	0x3E, 0x1B, 0x1F, 0x18, 0x25, 0x2F, 0x2C, 0x0A, 0x5D, 0x33, 0x07, 0x53,
	0x2A, 0x29, 0x71, 0x24, 0x4E, 0x14, 0x0E, 0x34, 0x28, 0x51, 0x37, 0x0F,
	0x38, 0x35, 0x17, 0x1B, 0x3E, 0x34, 0x09, 0x50, 0x2C, 0x08, 0x6D, 0x15,
	0x35, 0x14, 0x5C, 0x33, 0x5C, 0x4E, 0x06, 0x2C, 0x0B, 0x24, 0x0F, 0x2B,
	0x3E, 0x12, 0x3D, 0x32, 0x25, 0x24, 0x6D, 0x2B, 0x2A, 0x21, 0x21, 0x31,
	0x29, 0x38, 0x16, 0x28, 0x34, 0x38, 0x2C, 0x17, 0x22, 0x2F, 0x08, 0x52,
	0x45, 0x5A, 0x11, 0x3B, 0x0D, 0x5B, 0x59, 0x29, 0x1F, 0x59, 0x03, 0x27,
	0x0D, 0x2F, 0x59, 0x59, 0x1B, 0x11, 0x15, 0x08, 0x26, 0x40, 0x17, 0x47,
	0x34, 0x2D, 0x53, 0x3A, 0x1D, 0x4A, 0x0B, 0x1F, 0x25, 0x1E, 0x35, 0x08,
	0x27, 0x37, 0x5E, 0x16, 0x3D, 0x07, 0x27, 0x3A, 0x58, 0x16, 0x24, 0x2A,
	0x35, 0x54, 0x36, 0x3C, 0x7B, 0x21, 0x11, 0x23, 0x05, 0x74, 0x34, 0x2D,
	0x16, 0x18, 0x7B, 0x19, 0x0C, 0x3D, 0x04, 0x75, 0x1C, 0x14, 0x2F, 0x21,
	0x07, 0x1D, 0x24, 0x1F, 0x18, 0x77, 0x02, 0x36, 0x5E, 0x59, 0x0A, 0x03,
	0x09, 0x5E, 0x0D, 0x24, 0x3A, 0x2F, 0x04, 0x0F, 0x73, 0x0A, 0x0C, 0x16,
	0x26, 0x0A, 0x21, 0x00, 0x5E, 0x20, 0x36, 0x2E, 0x2D, 0x22, 0x0D, 0x3B,
	0x5B, 0x4E, 0x1C, 0x21, 0x33, 0x5D, 0x3B, 0x02, 0x13, 0x70, 0x1A, 0x07,
	0x16, 0x13, 0x03, 0x2D, 0x52, 0x1A, 0x13, 0x1B, 0x58, 0x24, 0x23, 0x3E,
	0x21, 0x54, 0x07, 0x1C, 0x20, 0x05, 0x5D, 0x19, 0x17, 0x2E, 0x2F, 0x3F,
	0x55, 0x27, 0x5B, 0x30, 0x2A, 0x00, 0x3D, 0x5D, 0x38, 0x2A, 0x10, 0x3C,
	0x24, 0x3B, 0x14, 0x02, 0x18, 0x3A, 0x2B, 0x43, 0x14, 0x2B, 0x09, 0x1A,
	0x58, 0x22, 0x58, 0x22, 0x14, 0x2F, 0x3B, 0x0F, 0x12, 0x34, 0x05, 0x39,
	0x3B, 0x0E, 0x09, 0x14, 0x32, 0x5A, 0x5A, 0x70, 0x09, 0x07, 0x5B, 0x32,
	0x25, 0x16, 0x50, 0x57, 0x1B, 0x3A, 0x39, 0x52, 0x5C, 0x3E, 0x31, 0x1B,
	0x33, 0x1C, 0x2C, 0x76, 0x27, 0x3B, 0x07, 0x3A, 0x73, 0x5D, 0x0F, 0x03,
	0x00, 0x00, 0x5C, 0x19, 0x2F, 0x3E, 0x05, 0x23, 0x08, 0x59, 0x23, 0x09,
	0x39, 0x56, 0x18, 0x2E, 0x26, 0x20, 0x4A, 0x45, 0x05, 0x73, 0x29, 0x0F,
	0x1B, 0x2D, 0x10, 0x23, 0x17, 0x20, 0x04, 0x03, 0x3B, 0x0F, 0x01, 0x5B,
	0x70, 0x39, 0x0E, 0x5A, 0x22, 0x0F, 0x07, 0x18, 0x38, 0x5A, 0x2E, 0x2B,
	0x59, 0x37, 0x26, 0x21, 0x06, 0x2F, 0x34, 0x03, 0x33, 0x3F, 0x55, 0x5A,
	0x19, 0x00, 0x5D, 0x19, 0x03, 0x38, 0x2D, 0x1A, 0x35, 0x01, 0x0A, 0x14,
	0x03, 0x11, 0x28, 0x2F, 0x2C, 0x15, 0x1B, 0x5E, 0x09, 0x20, 0x36, 0x2B,
	0x0A, 0x0A, 0x77, 0x15, 0x1B, 0x1E, 0x31, 0x27, 0x35, 0x51, 0x3B, 0x11,
	0x6D, 0x59, 0x12, 0x38, 0x13, 0x32, 0x04, 0x19, 0x57, 0x1D, 0x16, 0x55,
	0x2A, 0x57, 0x20, 0x07, 0x35, 0x2C, 0x23, 0x32, 0x25, 0x0D, 0x00, 0x0D,
	0x3A, 0x70, 0x22, 0x25, 0x57, 0x40, 0x33, 0x02, 0x27, 0x09, 0x53, 0x20,
	0x35, 0x02, 0x0A, 0x18, 0x1B, 0x5A, 0x25, 0x2A, 0x1C, 0x0C, 0x1C, 0x2F,
	0x1E, 0x2C, 0x24, 0x06, 0x2E, 0x09, 0x33, 0x37, 0x03, 0x17, 0x22, 0x2C,
	0x14, 0x20, 0x1B, 0x56, 0x2C, 0x29, 0x21, 0x15, 0x21, 0x0C, 0x7B, 0x35,
	0x2F, 0x17, 0x24, 0x38, 0x29, 0x58, 0x58, 0x5B, 0x11, 0x05, 0x50, 0x17,
	0x3F, 0x32, 0x38, 0x20, 0x08, 0x38, 0x36, 0x1B, 0x27, 0x58, 0x1C, 0x25,
	0x1B, 0x4E, 0x17, 0x28, 0x18, 0x5E, 0x05, 0x3D, 0x19, 0x18, 0x19, 0x33,
	0x24, 0x3D, 0x28, 0x38, 0x36, 0x58, 0x13, 0x20, 0x1F, 0x2F, 0x29, 0x20,
	0x33, 0x27, 0x05, 0x1D, 0x13, 0x20, 0x2D, 0x36, 0x45, 0x3E, 0x10, 0x5C,
	0x2F, 0x18, 0x3E, 0x30, 0x03, 0x4A, 0x3D, 0x00, 0x0B, 0x1D, 0x17, 0x05,
	0x03, 0x35, 0x08, 0x02, 0x0C, 0x33, 0x33, 0x22, 0x0B, 0x37, 0x20, 0x09,
	0x5D, 0x51, 0x24, 0x05, 0x10, 0x18, 0x0F, 0x05, 0x32, 0x20, 0x47, 0x53,
	0x3D, 0x19, 0x1A, 0x1B, 0x19, 0x23, 0x5C, 0x14, 0x5E, 0x58, 0x27, 0x3B,
	0x25, 0x5F, 0x1B, 0x1B, 0x27, 0x00, 0x1B, 0x20, 0x2B, 0x1C, 0x26, 0x06,
	0x18, 0x0C, 0x2A, 0x14, 0x26, 0x16, 0x5C, 0x3A, 0x21, 0x5A, 0x2D, 0x06,
	0x28, 0x33, 0x3D, 0x11, 0x45, 0x3C, 0x26, 0x3E, 0x2D, 0x06, 0x44, 0x72,
	0x22, 0x18, 0x02, 0x2C, 0x34, 0x0B, 0x05, 0x58, 0x3D, 0x04, 0x18, 0x12,
	0x16, 0x25, 0x13, 0x20, 0x26, 0x2C, 0x0C, 0x0C, 0x5B, 0x07, 0x01, 0x44,
	0x26, 0x5C, 0x06, 0x36, 0x19, 0x08, 0x1E, 0x52, 0x1E, 0x28, 0x28, 0x08,
	0x38, 0x34, 0x3C, 0x27, 0x3D, 0x57, 0x1A, 0x52, 0x14, 0x1D, 0x30, 0x20,
	0x24, 0x1B, 0x04, 0x16, 0x38, 0x1A, 0x2E, 0x38, 0x1B, 0x3F, 0x5A, 0x20,
	0x0A, 0x1B, 0x38, 0x53, 0x13, 0x59, 0x0A, 0x0A, 0x08, 0x01, 0x59, 0x2A,
	0x00, 0x0A, 0x01, 0x18, 0x2E, 0x57, 0x1B, 0x38, 0x06, 0x18, 0x57, 0x44,
	0x03, 0x5A, 0x09, 0x2B, 0x2D, 0x0F, 0x5B, 0x13, 0x08, 0x0F, 0x10, 0x0E,
	0x59, 0x34, 0x38, 0x75, 0x54, 0x15, 0x38, 0x02, 0x26, 0x27, 0x18, 0x45,
	0x5A, 0x2A, 0x54, 0x17, 0x1E, 0x26, 0x7B, 0x58, 0x4E, 0x5E, 0x59, 0x7A,
	0x2F, 0x15, 0x3B, 0x0A, 0x03, 0x3E, 0x33, 0x27, 0x2F, 0x12, 0x2B, 0x4A,
	0x58, 0x1C, 0x1A, 0x3F, 0x00, 0x2C, 0x5C, 0x27, 0x06, 0x06, 0x02, 0x1D,
	0x26, 0x34, 0x02, 0x1E, 0x3B, 0x09, 0x3E, 0x36, 0x02, 0x38, 0x0D, 0x3A,
	0x54, 0x57, 0x11, 0x25, 0x2A, 0x4E, 0x5D, 0x20, 0x00, 0x28, 0x16, 0x21,
	0x03, 0x0D, 0x27, 0x55, 0x18, 0x58, 0x2F, 0x27, 0x14, 0x22, 0x1A, 0x04,
	0x36, 0x05, 0x59, 0x2D, 0x73, 0x28, 0x30, 0x21, 0x32, 0x03, 0x2B, 0x38,
	0x0B, 0x0D, 0x26, 0x5D, 0x29, 0x25, 0x25, 0x21, 0x04, 0x2B, 0x02, 0x58,
	0x00, 0x3A, 0x07, 0x22, 0x29, 0x0A, 0x59, 0x2F, 0x18, 0x29, 0x0A, 0x5F,
	0x22, 0x5D, 0x0F, 0x11, 0x59, 0x0D, 0x5C, 0x39, 0x71, 0x55, 0x28, 0x5A,
	0x3A, 0x17, 0x06, 0x52, 0x37, 0x1C, 0x75, 0x0F, 0x4E, 0x37, 0x5A, 0x2D,
	0x58, 0x2F, 0x00, 0x0D, 0x0B, 0x2A, 0x11, 0x25, 0x0E, 0x1B, 0x47, 0x22,
	0x29, 0x5B, 0x77, 0x0E, 0x05, 0x27, 0x11, 0x03, 0x07, 0x1B, 0x22, 0x29,
	0x06, 0x20, 0x12, 0x5E, 0x38, 0x18, 0x3E, 0x2D, 0x02, 0x58, 0x7B, 0x59,
	0x20, 0x27, 0x1B, 0x00, 0x3E, 0x2F, 0x06, 0x5B, 0x24, 0x1D, 0x1B, 0x29,
	0x01, 0x29, 0x09, 0x0B, 0x23, 0x0D, 0x24, 0x19, 0x32, 0x0D, 0x22, 0x26,
	0x0D, 0x33, 0x56, 0x3E, 0x71, 0x05, 0x0F, 0x1D, 0x1A, 0x3A, 0x35, 0x15,
	0x1B, 0x5E, 0x1B, 0x5D, 0x2C, 0x2C, 0x3B, 0x00, 0x3E, 0x58, 0x26, 0x5D,
	0x69, 0x3A, 0x50, 0x1C, 0x3E, 0x11, 0x0F, 0x29, 0x25, 0x11, 0x01, 0x01,
	0x2D, 0x06, 0x0F, 0x29, 0x29, 0x4E, 0x45, 0x31, 0x34, 0x05, 0x13, 0x0C,
	0x03, 0x7B, 0x0E, 0x22, 0x08, 0x26, 0x20, 0x35, 0x52, 0x0D, 0x5B, 0x0D,
	0x5F, 0x0D, 0x5A, 0x33, 0x07, 0x00, 0x1B, 0x0A, 0x3E, 0x24, 0x43, 0x17,
	0x2D, 0x20, 0x75, 0x0E, 0x14, 0x3E, 0x2A, 0x73, 0x47, 0x52, 0x14, 0x32,
	0x2F, 0x1F, 0x50, 0x59, 0x08, 0x2A, 0x2B, 0x32, 0x0D, 0x01, 0x76, 0x19,
	0x50, 0x19, 0x0D, 0x36, 0x19, 0x27, 0x5A, 0x58, 0x1B, 0x5A, 0x34, 0x34,
	0x09, 0x0E, 0x5E, 0x4A, 0x03, 0x24, 0x0F, 0x1F, 0x23, 0x3D, 0x2E, 0x2A,
	0x43, 0x3B, 0x22, 0x12, 0x74, 0x1C, 0x32, 0x09, 0x5E, 0x03, 0x03, 0x32,
	0x07, 0x08, 0x0D, 0x59, 0x23, 0x58, 0x33, 0x15, 0x26, 0x28, 0x59, 0x5E,
	0x18, 0x55, 0x14, 0x01, 0x2F, 0x2A, 0x26, 0x00, 0x0A, 0x5A, 0x37, 0x00,
	0x2E, 0x1E, 0x39, 0x21, 0x24, 0x22, 0x07, 0x31, 0x0C, 0x06, 0x0F, 0x01,
	0x26, 0x12, 0x1B, 0x0B, 0x3B, 0x5E, 0x28, 0x3D, 0x0C, 0x09, 0x2D, 0x11,
	0x06, 0x34, 0x3E, 0x5D, 0x04, 0x00, 0x54, 0x16, 0x13, 0x77, 0x38, 0x12,
	0x25, 0x09, 0x10, 0x3A, 0x30, 0x5D, 0x0A, 0x15, 0x2F, 0x32, 0x2D, 0x11,
	0x0E, 0x1C, 0x0C, 0x07, 0x12, 0x74, 0x16, 0x54, 0x2D, 0x11, 0x06, 0x05,
	0x39, 0x14, 0x07, 0x3B, 0x27, 0x58, 0x0A, 0x2A, 0x70, 0x1C, 0x2C, 0x06,
	0x08, 0x24, 0x3A, 0x31, 0x00, 0x28, 0x23, 0x19, 0x31, 0x06, 0x3D, 0x0C,
	0x1E, 0x39, 0x1C, 0x40, 0x05, 0x25, 0x37, 0x1F, 0x1C, 0x03, 0x0B, 0x34,
	0x3B, 0x2F, 0x14, 0x04, 0x2B, 0x08, 0x52, 0x37, 0x0F, 0x17, 0x0F, 0x5F,
	0x17, 0x5F, 0x0E, 0x0B, 0x0A, 0x0D, 0x5F, 0x54, 0x26, 0x5E, 0x0E, 0x5B,
	0x2C, 0x2C, 0x2F, 0x0E, 0x5B, 0x35, 0x41, 0x09, 0x0A, 0x2E, 0x2D, 0x59,
	0x38, 0x30, 0x3A, 0x38, 0x14, 0x19, 0x21, 0x3C, 0x53, 0x16, 0x1B, 0x29,
	0x58, 0x28, 0x56, 0x26, 0x35, 0x00, 0x25, 0x21, 0x24, 0x38, 0x38, 0x56,
	0x2A, 0x08, 0x25, 0x2B, 0x20, 0x2C, 0x3B, 0x32, 0x2E, 0x26, 0x3E, 0x01,
	0x7B, 0x1E, 0x14, 0x24, 0x01, 0x1B, 0x18, 0x02, 0x2C, 0x3C, 0x12, 0x06,
	0x10, 0x5E, 0x21, 0x69, 0x5F, 0x1B, 0x2C, 0x18, 0x10, 0x5F, 0x22, 0x34,
	0x40, 0x36, 0x0E, 0x26, 0x00, 0x32, 0x26, 0x2E, 0x2A, 0x14, 0x07, 0x71,
	0x04, 0x59, 0x1A, 0x5C, 0x25, 0x3F, 0x57, 0x25, 0x2E, 0x2E, 0x3A, 0x18,
	0x02, 0x08, 0x13, 0x55, 0x24, 0x18, 0x32, 0x00, 0x08, 0x15, 0x19, 0x13,
	0x0E, 0x28, 0x0A, 0x29, 0x38, 0x33, 0x1E, 0x29, 0x09, 0x1D, 0x23, 0x03,
	0x0A, 0x20, 0x27, 0x3A, 0x21, 0x17, 0x1F, 0x21, 0x0F, 0x01, 0x0A, 0x04,
	0x33, 0x77, 0x0F, 0x53, 0x2A, 0x07, 0x33, 0x28, 0x55, 0x05, 0x32, 0x05,
	0x29, 0x1B, 0x0D, 0x1E, 0x31, 0x0B, 0x26, 0x1F, 0x0F, 0x70, 0x18, 0x51,
	0x1F, 0x5D, 0x29, 0x1C, 0x32, 0x5B, 0x06, 0x23, 0x5C, 0x0F, 0x5C, 0x3C,
	0x31, 0x3F, 0x3B, 0x5F, 0x3E, 0x04, 0x09, 0x38, 0x08, 0x2C, 0x2B, 0x34,
	0x00, 0x06, 0x13, 0x76, 0x2D, 0x23, 0x17, 0x01, 0x36, 0x0A, 0x08, 0x45,
	0x02, 0x08, 0x3D, 0x31, 0x3D, 0x5A, 0x29, 0x07, 0x4E, 0x27, 0x1A, 0x25,
	0x0A, 0x28, 0x04, 0x05, 0x2C, 0x5A, 0x52, 0x3D, 0x0F, 0x69, 0x1D, 0x51,
	0x1D, 0x2F, 0x3B, 0x15, 0x14, 0x29, 0x3A, 0x74, 0x59, 0x2E, 0x05, 0x00,
	0x1A, 0x1B, 0x0D, 0x3D, 0x01, 0x04, 0x3D, 0x0F, 0x01, 0x05, 0x35, 0x00,
	0x32, 0x26, 0x00, 0x3A, 0x20, 0x32, 0x07, 0x0A, 0x32, 0x43, 0x17, 0x2B,
	0x08, 0x12, 0x02, 0x10, 0x14, 0x1A, 0x77, 0x1B, 0x4A, 0x3D, 0x04, 0x2C,
	0x34, 0x2D, 0x5A, 0x0A, 0x73, 0x07, 0x39, 0x5C, 0x2E, 0x23, 0x25, 0x00,
	0x25, 0x52, 0x2F, 0x07, 0x06, 0x24, 0x5D, 0x70, 0x0E, 0x34, 0x0C, 0x29,
	0x36, 0x59, 0x13, 0x5D, 0x07, 0x05, 0x26, 0x06, 0x0C, 0x12, 0x03, 0x05,
	0x04, 0x08, 0x02, 0x15, 0x16, 0x34, 0x3C, 0x02, 0x75, 0x47, 0x23, 0x1D,
	0x09, 0x29, 0x24, 0x56, 0x28, 0x39, 0x09, 0x3B, 0x4A, 0x00, 0x5F, 0x0A,
	0x2B, 0x56, 0x57, 0x06, 0x2E, 0x22, 0x14, 0x24, 0x01, 0x28, 0x5C, 0x50,
	0x0B, 0x5A, 0x2A, 0x07, 0x09, 0x03, 0x11, 0x72, 0x3D, 0x2A, 0x28, 0x2E,
	0x10, 0x3C, 0x25, 0x3B, 0x27, 0x33, 0x07, 0x38, 0x0C, 0x2E, 0x36, 0x14,
	0x15, 0x38, 0x1C, 0x38, 0x3B, 0x2C, 0x39, 0x26, 0x03, 0x1F, 0x12, 0x56,
	0x07, 0x12, 0x23, 0x22, 0x41, 0x27, 0x09, 0x0E, 0x19, 0x22, 0x18, 0x07,
	0x09, 0x04, 0x2D, 0x06, 0x28, 0x04, 0x25, 0x41, 0x31, 0x00, 0x1D, 0x2F,
	0x20, 0x11, 0x2A, 0x43, 0x11, 0x28, 0x0C, 0x14, 0x14, 0x57, 0x2C, 0x0E,
	0x77, 0x39, 0x3B, 0x18, 0x2D, 0x23, 0x02, 0x2E, 0x17, 0x06, 0x13, 0x24,
	0x20, 0x2B, 0x02, 0x1A, 0x01, 0x15, 0x3B, 0x31, 0x70, 0x06, 0x4E, 0x1B,
	0x2E, 0x15, 0x47, 0x32, 0x24, 0x53, 0x04, 0x0F, 0x55, 0x06, 0x2E, 0x37,
	0x2A, 0x26, 0x45, 0x12, 0x26, 0x2F, 0x33, 0x57, 0x32, 0x18, 0x21, 0x04,
	0x0D, 0x25, 0x35, 0x01, 0x54, 0x0F, 0x3D, 0x2F, 0x2E, 0x2B, 0x22, 0x44,
	0x2E, 0x35, 0x23, 0x2D, 0x2F, 0x32, 0x3F, 0x16, 0x01, 0x3D, 0x7A, 0x22,
	0x30, 0x5F, 0x19, 0x15, 0x24, 0x55, 0x1E, 0x53, 0x07, 0x0F, 0x33, 0x0C,
	0x1A, 0x2D, 0x3B, 0x4A, 0x3B, 0x3D, 0x35, 0x38, 0x34, 0x34, 0x20, 0x07,
	0x27, 0x4E, 0x1F, 0x24, 0x25, 0x1C, 0x2F, 0x36, 0x32, 0x0A, 0x28, 0x18,
	0x3E, 0x0E, 0x13, 0x2A, 0x06, 0x22, 0x24, 0x0B, 0x07, 0x53, 0x0A, 0x2D,
	0x35, 0x3D, 0x04, 0x58, 0x59, 0x33, 0x24, 0x2A, 0x26, 0x38, 0x3B, 0x03,
	0x4A, 0x25, 0x29, 0x0B, 0x0B, 0x00, 0x39, 0x5C, 0x12, 0x5A, 0x20, 0x20,
	0x11, 0x73, 0x0A, 0x17, 0x1A, 0x1D, 0x07, 0x0E, 0x0E, 0x5C, 0x28, 0x36,
	0x08, 0x0F, 0x38, 0x2D, 0x35, 0x38, 0x2A, 0x2C, 0x1B, 0x1B, 0x1C, 0x00,
	0x3F, 0x23, 0x2E, 0x0F, 0x0B, 0x5E, 0x19, 0x72, 0x05, 0x57, 0x09, 0x53,
	0x34, 0x1D, 0x2A, 0x1E, 0x5D, 0x18, 0x2B, 0x03, 0x1D, 0x05, 0x2A, 0x14,
	0x08, 0x5D, 0x5C, 0x3A, 0x29, 0x55, 0x23, 0x1E, 0x31, 0x3B, 0x03, 0x58,
	0x1F, 0x2F, 0x18, 0x32, 0x07, 0x06, 0x1B, 0x26, 0x12, 0x09, 0x2A, 0x6D,
	0x20, 0x0C, 0x01, 0x09, 0x35, 0x5B, 0x15, 0x26, 0x39, 0x33, 0x2A, 0x0A,
	0x20, 0x27, 0x17, 0x2B, 0x10, 0x1B, 0x44, 0x0E, 0x1E, 0x51, 0x26, 0x44,
	0x2F, 0x2E, 0x16, 0x39, 0x39, 0x71, 0x25, 0x10, 0x0F, 0x2A, 0x04, 0x01,
	0x00, 0x3D, 0x0E, 0x27, 0x2F, 0x55, 0x5D, 0x06, 0x0F, 0x2F, 0x0E, 0x2D,
	0x0A, 0x03, 0x23, 0x36, 0x09, 0x5F, 0x17, 0x3C, 0x38, 0x37, 0x01, 0x00,
	0x03, 0x13, 0x0F, 0x13, 0x00, 0x34, 0x54, 0x1E, 0x1B, 0x70, 0x36, 0x0F,
	0x21, 0x03, 0x09, 0x5E, 0x4E, 0x41, 0x31, 0x06, 0x1A, 0x07, 0x28, 0x08,
	0x76, 0x08, 0x04, 0x06, 0x38, 0x1A, 0x3A, 0x56, 0x1B, 0x27, 0x3A, 0x0D,
	0x0F, 0x38, 0x07, 0x0E, 0x54, 0x13, 0x21, 0x11, 0x27, 0x01, 0x10, 0x28,
	0x27, 0x21, 0x5A, 0x2C, 0x3F, 0x13, 0x71, 0x20, 0x14, 0x5F, 0x40, 0x0E,
	0x03, 0x09, 0x04, 0x0C, 0x10, 0x3F, 0x50, 0x04, 0x2C, 0x03, 0x20, 0x1B,
	0x29, 0x58, 0x3A, 0x0F, 0x2A, 0x3B, 0x0A, 0x04, 0x19, 0x34, 0x04, 0x3C,
	0x2F, 0x18, 0x2D, 0x5E, 0x0C, 0x3B, 0x2E, 0x00, 0x09, 0x44, 0x25, 0x14,
	0x28, 0x18, 0x24, 0x09, 0x06, 0x08, 0x0B, 0x2F, 0x77, 0x20, 0x08, 0x20,
	0x2A, 0x2F, 0x05, 0x58, 0x0D, 0x1D, 0x75, 0x21, 0x26, 0x1D, 0x2D, 0x11,
	0x04, 0x4E, 0x0F, 0x07, 0x35, 0x07, 0x0B, 0x59, 0x00, 0x2F, 0x54, 0x06,
	0x07, 0x1F, 0x03, 0x3A, 0x11, 0x2D, 0x00, 0x70, 0x0F, 0x05, 0x5D, 0x18,
	0x11, 0x14, 0x02, 0x5F, 0x40, 0x73, 0x27, 0x35, 0x2C, 0x3D, 0x24, 0x1A,
	0x35, 0x01, 0x5E, 0x71, 0x36, 0x18, 0x24, 0x5A, 0x14, 0x1F, 0x32, 0x23,
	0x2D, 0x27, 0x34, 0x3B, 0x26, 0x2C, 0x15, 0x25, 0x12, 0x22, 0x04, 0x74,
	0x3D, 0x29, 0x0A, 0x26, 0x10, 0x47, 0x02, 0x5E, 0x5B, 0x09, 0x34, 0x2C,
	0x1F, 0x2E, 0x37, 0x55, 0x24, 0x0F, 0x33, 0x18, 0x54, 0x15, 0x2D, 0x02,
	0x0C, 0x20, 0x2D, 0x1E, 0x1B, 0x34, 0x3B, 0x04, 0x25, 0x12, 0x34, 0x2B,
	0x59, 0x5B, 0x5E, 0x1A, 0x3F, 0x24, 0x21, 0x19, 0x26, 0x36, 0x36, 0x06,
	0x0A, 0x28, 0x36, 0x55, 0x26, 0x22, 0x0E, 0x3C, 0x05, 0x3C, 0x5F, 0x0C,
	0x3F, 0x0A, 0x05, 0x2C, 0x26, 0x5E, 0x52, 0x45, 0x08, 0x05, 0x28, 0x0C,
	0x38, 0x03, 0x10, 0x25, 0x56, 0x1B, 0x26, 0x31, 0x00, 0x38, 0x39, 0x5C,
	0x7A, 0x0D, 0x53, 0x5E, 0x33, 0x71, 0x18, 0x3B, 0x0D, 0x2A, 0x32, 0x1D,
	0x14, 0x28, 0x5E, 0x35, 0x3A, 0x0A, 0x2F, 0x31, 0x27, 0x0A, 0x55, 0x27,
	0x58, 0x1B, 0x1C, 0x51, 0x05, 0x0A, 0x3A, 0x25, 0x02, 0x17, 0x13, 0x1B,
	0x0E, 0x3B, 0x05, 0x22, 0x13, 0x1C, 0x4A, 0x1C, 0x05, 0x21, 0x19, 0x31,
	0x1D, 0x13, 0x23, 0x18, 0x0B, 0x2F, 0x06, 0x0F, 0x58, 0x58, 0x5F, 0x44,
	0x73, 0x5C, 0x51, 0x09, 0x0F, 0x74, 0x22, 0x04, 0x58, 0x1C, 0x10, 0x07,
	0x17, 0x5B, 0x2F, 0x06, 0x34, 0x36, 0x5F, 0x20, 0x2D, 0x3C, 0x2C, 0x2B,
	0x3B, 0x29, 0x5B, 0x24, 0x1C, 0x2C, 0x70, 0x06, 0x02, 0x21, 0x05, 0x09,
	0x2B, 0x0D, 0x0A, 0x1C, 0x34, 0x03, 0x2D, 0x2A, 0x5F, 0x0E, 0x01, 0x59,
	0x0B, 0x12, 0x08, 0x5C, 0x39, 0x3A, 0x1D, 0x0B, 0x59, 0x11, 0x2F, 0x20,
	0x06, 0x22, 0x28, 0x04, 0x18, 0x1B, 0x27, 0x0A, 0x36, 0x23, 0x0C, 0x0D,
	0x27, 0x2D, 0x0E, 0x23, 0x2B, 0x2E, 0x27, 0x2D, 0x18, 0x1F, 0x59, 0x1B,
	0x0A, 0x2A, 0x1A, 0x29, 0x0B, 0x40, 0x23, 0x05, 0x38, 0x39, 0x3A, 0x04,
	0x2B, 0x05, 0x58, 0x00, 0x2C, 0x0E, 0x18, 0x1A, 0x39, 0x26, 0x5F, 0x07,
	0x29, 0x09, 0x0E, 0x43, 0x39, 0x19, 0x38, 0x14, 0x2E, 0x30, 0x26, 0x07,
	0x69, 0x35, 0x0E, 0x28, 0x0D, 0x01, 0x16, 0x54, 0x07, 0x04, 0x00, 0x3E,
	0x09, 0x09, 0x2A, 0x03, 0x2B, 0x32, 0x1A, 0x2F, 0x2C, 0x1F, 0x38, 0x2C,
	0x33, 0x07, 0x28, 0x4A, 0x3F, 0x40, 0x29, 0x3F, 0x1B, 0x59, 0x32, 0x3A,
	0x43, 0x2A, 0x2B, 0x28, 0x0F, 0x24, 0x50, 0x3B, 0x13, 0x2C, 0x23, 0x27,
	0x58, 0x0A, 0x31, 0x29, 0x55, 0x5F, 0x33, 0x1B, 0x5E, 0x0B, 0x3C, 0x02,
	0x35, 0x2B, 0x38, 0x5E, 0x5A, 0x1B, 0x2F, 0x18, 0x0B, 0x02, 0x2A, 0x07,
	0x13, 0x17, 0x11, 0x0D, 0x05, 0x59, 0x2B, 0x3F, 0x2B, 0x28, 0x09, 0x21,
	0x40, 0x0B, 0x26, 0x25, 0x36, 0x09, 0x14, 0x26, 0x4E, 0x3D, 0x19, 0x0B,
	0x3C, 0x57, 0x3A, 0x52, 0x23, 0x05, 0x24, 0x0B, 0x27, 0x74, 0x2D, 0x3B,
	0x26, 0x32, 0x35, 0x01, 0x24, 0x56, 0x3B, 0x6D, 0x35, 0x04, 0x56, 0x52,
	0x2D, 0x27, 0x2D, 0x0F, 0x1E, 0x21, 0x0A, 0x33, 0x0D, 0x13, 0x2B, 0x2B,
	0x25, 0x05, 0x25, 0x14, 0x1F, 0x2C, 0x2D, 0x04, 0x2D, 0x27, 0x25, 0x3D,
	0x24, 0x35, 0x1E, 0x32, 0x2C, 0x0C, 0x1B, 0x08, 0x08, 0x02, 0x39, 0x10,
	0x2A, 0x20, 0x37, 0x32, 0x2B, 0x1F, 0x20, 0x23, 0x3F, 0x33, 0x29, 0x0E,
	0x27, 0x2A, 0x33, 0x03, 0x55, 0x19, 0x03, 0x2B, 0x5B, 0x4E, 0x5D, 0x0A,
	0x27, 0x54, 0x02, 0x1B, 0x3C, 0x0F, 0x2E, 0x18, 0x28, 0x3D, 0x07, 0x3E,
	0x2E, 0x41, 0x31, 0x00, 0x1A, 0x31, 0x0F, 0x28, 0x28, 0x0A, 0x0A, 0x00,
	0x24, 0x15, 0x09, 0x26, 0x0D, 0x1F, 0x1A, 0x1A, 0x04, 0x59, 0x40, 0x71,
	0x5D, 0x0D, 0x1A, 0x1D, 0x34, 0x0A, 0x04, 0x0C, 0x39, 0x26, 0x04, 0x2B,
	0x3A, 0x00, 0x74, 0x15, 0x12, 0x59, 0x24, 0x38, 0x1F, 0x54, 0x21, 0x3F,
	0x75, 0x2A, 0x09, 0x2A, 0x06, 0x7B, 0x03, 0x05, 0x2A, 0x3D, 0x30, 0x3B,
	0x06, 0x07, 0x00, 0x23, 0x3A, 0x2D, 0x3D, 0x2E, 0x35, 0x23, 0x55, 0x56,
	0x09, 0x25, 0x23, 0x2A, 0x2F, 0x0A, 0x72, 0x29, 0x0A, 0x3F, 0x23, 0x17,
	0x0E, 0x57, 0x02, 0x1F, 0x08, 0x54, 0x02, 0x00, 0x0A, 0x0A, 0x28, 0x56,
	0x21, 0x21, 0x33, 0x05, 0x02, 0x39, 0x2C, 0x26, 0x27, 0x54, 0x2B, 0x07,
	0x3B, 0x5F, 0x03, 0x27, 0x33, 0x24, 0x1D, 0x00, 0x1E, 0x2A, 0x71, 0x1C,
	0x2E, 0x41, 0x2A, 0x35, 0x16, 0x0A, 0x1E, 0x33, 0x17, 0x20, 0x3B, 0x27,
	0x01, 0x16, 0x2D, 0x0B, 0x14, 0x31, 0x03, 0x38, 0x14, 0x03, 0x3C, 0x18,
	0x25, 0x11, 0x56, 0x11, 0x69, 0x24, 0x0A, 0x0D, 0x01, 0x27, 0x03, 0x06,
	0x57, 0x44, 0x11, 0x23, 0x56, 0x16, 0x19, 0x04, 0x5F, 0x1B, 0x07, 0x02,
	0x35, 0x34, 0x23, 0x04, 0x08, 0x73, 0x25, 0x2F, 0x58, 0x23, 0x71, 0x27,
	0x0D, 0x24, 0x32, 0x2C, 0x3C, 0x4A, 0x3F, 0x11, 0x35, 0x0F, 0x4E, 0x05,
	0x3F, 0x12, 0x2D, 0x13, 0x2A, 0x09, 0x04, 0x14, 0x08, 0x45, 0x0F, 0x12,
	0x36, 0x31, 0x28, 0x20, 0x36, 0x04, 0x58, 0x2A, 0x39, 0x17, 0x2E, 0x56,
	0x34, 0x2A, 0x27, 0x3E, 0x37, 0x58, 0x58, 0x04, 0x0B, 0x32, 0x2D, 0x52,
	0x69, 0x2D, 0x22, 0x5E, 0x02, 0x12, 0x1E, 0x55, 0x34, 0x5D, 0x24, 0x14,
	0x22, 0x38, 0x3E, 0x17, 0x3A, 0x33, 0x58, 0x3A, 0x36, 0x1F, 0x16, 0x26,
	0x3B, 0x33, 0x55, 0x23, 0x2C, 0x1A, 0x74, 0x1E, 0x18, 0x39, 0x32, 0x30,
	0x04, 0x05, 0x0B, 0x21, 0x29, 0x23, 0x30, 0x3F, 0x2C, 0x2D, 0x2F, 0x54,
	0x34, 0x2D, 0x6D, 0x58, 0x0C, 0x29, 0x2A, 0x74, 0x36, 0x22, 0x0D, 0x38,
	0x10, 0x2A, 0x39, 0x2D, 0x19, 0x24, 0x1A, 0x58, 0x2B, 0x13, 0x1A, 0x1C,
	0x00, 0x29, 0x33, 0x35, 0x27, 0x24, 0x2A, 0x27, 0x26, 0x2E, 0x23, 0x20,
	0x02, 0x06, 0x29, 0x56, 0x03, 0x03, 0x17, 0x5C, 0x04, 0x2D, 0x1A, 0x69,
	0x1D, 0x0B, 0x09, 0x1F, 0x27, 0x0B, 0x00, 0x3D, 0x5D, 0x0B, 0x5C, 0x57,
	0x22, 0x20, 0x29, 0x2B, 0x25, 0x1A, 0x5B, 0x71, 0x39, 0x2A, 0x23, 0x38,
	0x73, 0x14, 0x08, 0x45, 0x2A, 0x71, 0x58, 0x19, 0x5D, 0x28, 0x34, 0x1F,
	0x17, 0x21, 0x18, 0x03, 0x3E, 0x0D, 0x16, 0x01, 0x27, 0x26, 0x04, 0x5A,
	0x44, 0x36, 0x1C, 0x57, 0x5B, 0x1C, 0x05, 0x5C, 0x23, 0x0D, 0x3F, 0x2B,
	0x58, 0x20, 0x2B, 0x26, 0x1A, 0x34, 0x58, 0x0A, 0x40, 0x1B, 0x24, 0x26,
	0x23, 0x5A, 0x16, 0x1C, 0x05, 0x26, 0x58, 0x2A, 0x09, 0x04, 0x2F, 0x1E,
	0x32, 0x55, 0x22, 0x0F, 0x11, 0x2C, 0x3B, 0x4E, 0x38, 0x31, 0x01, 0x01,
	0x11, 0x58, 0x1C, 0x29, 0x1A, 0x4E, 0x59, 0x5D, 0x0B, 0x1E, 0x1B, 0x23,
	0x28, 0x73, 0x59, 0x4E, 0x08, 0x32, 0x18, 0x3B, 0x36, 0x01, 0x5C, 0x05,
	0x5F, 0x22, 0x37, 0x0D, 0x33, 0x16, 0x11, 0x29, 0x24, 0x10, 0x3C, 0x16,
	0x16, 0x3D, 0x24, 0x15, 0x4E, 0x05, 0x27, 0x0A, 0x2D, 0x4E, 0x2C, 0x12,
	0x3A, 0x2F, 0x2B, 0x2A, 0x23, 0x1A, 0x04, 0x58, 0x01, 0x3A, 0x31, 0x3E,
	0x51, 0x3E, 0x31, 0x01, 0x14, 0x07, 0x41, 0x05, 0x70, 0x5A, 0x59, 0x5F,
	0x44, 0x0F, 0x34, 0x37, 0x5B, 0x24, 0x71, 0x34, 0x1B, 0x0B, 0x39, 0x36,
	0x59, 0x57, 0x17, 0x00, 0x72, 0x55, 0x22, 0x01, 0x07, 0x17, 0x1E, 0x52,
	0x1F, 0x5D, 0x04, 0x55, 0x3B, 0x5C, 0x07, 0x00, 0x1F, 0x59, 0x14, 0x1E,
	0x2E, 0x5E, 0x06, 0x38, 0x13, 0x05, 0x5F, 0x0F, 0x56, 0x21, 0x08, 0x1C,
	0x3B, 0x3C, 0x5A, 0x05, 0x09, 0x05, 0x09, 0x0A, 0x25, 0x2E, 0x23, 0x25,
	0x13, 0x33, 0x28, 0x54, 0x3F, 0x02, 0x37, 0x09, 0x26, 0x18, 0x2F, 0x37,
	0x0D, 0x54, 0x2C, 0x18, 0x74, 0x5F, 0x58, 0x23, 0x39, 0x2C, 0x2B, 0x4E,
	0x22, 0x09, 0x6D, 0x18, 0x4E, 0x2B, 0x44, 0x08, 0x00, 0x2F, 0x5F, 0x1D,
	0x35, 0x55, 0x17, 0x21, 0x44, 0x77, 0x3F, 0x24, 0x58, 0x05, 0x74, 0x1C,
	0x00, 0x3E, 0x01, 0x34, 0x07, 0x10, 0x2C, 0x5C, 0x30, 0x59, 0x34, 0x5F,
	0x58, 0x0F, 0x54, 0x34, 0x03, 0x3E, 0x00, 0x1E, 0x12, 0x59, 0x29, 0x37,
	0x34, 0x00, 0x57, 0x20, 0x00, 0x2A, 0x34, 0x2A, 0x05, 0x0A, 0x26, 0x04,
	0x39, 0x3A, 0x29, 0x09, 0x32, 0x06, 0x3F, 0x23, 0x5D, 0x06, 0x0F, 0x38,
	0x3A, 0x5E, 0x33, 0x2C, 0x1B, 0x69, 0x0B, 0x11, 0x04, 0x07, 0x27, 0x06,
	0x36, 0x3B, 0x20, 0x2F, 0x27, 0x25, 0x02, 0x19, 0x00, 0x5B, 0x07, 0x26,
	0x1C, 0x75, 0x1F, 0x0D, 0x39, 0x0C, 0x10, 0x25, 0x06, 0x3B, 0x25, 0x34,
	0x18, 0x27, 0x58, 0x3F, 0x73, 0x1F, 0x07, 0x41, 0x40, 0x71, 0x14, 0x11,
	0x5F, 0x5C, 0x70, 0x02, 0x50, 0x1B, 0x19, 0x33, 0x39, 0x2A, 0x0B, 0x53,
	0x38, 0x29, 0x1B, 0x58, 0x03, 0x2D, 0x35, 0x53, 0x1A, 0x22, 0x23, 0x5F,
	0x25, 0x29, 0x1A, 0x20, 0x22, 0x4E, 0x5D, 0x27, 0x27, 0x38, 0x0B, 0x56,
	0x00, 0x32, 0x1C, 0x51, 0x36, 0x5C, 0x30, 0x24, 0x24, 0x37, 0x13, 0x7A,
	0x3F, 0x08, 0x09, 0x3C, 0x26, 0x1F, 0x37, 0x5F, 0x01, 0x2F, 0x05, 0x13,
	0x06, 0x5C, 0x13, 0x0A, 0x23, 0x36, 0x3D, 0x13, 0x00, 0x17, 0x09, 0x13,
	0x23, 0x3D, 0x32, 0x1D, 0x11, 0x10, 0x2A, 0x10, 0x19, 0x3D, 0x76, 0x0D,
	0x38, 0x2A, 0x32, 0x70, 0x5D, 0x00, 0x14, 0x01, 0x2A, 0x0F, 0x57, 0x0C,
	0x24, 0x04, 0x19, 0x32, 0x26, 0x3A, 0x29, 0x54, 0x08, 0x22, 0x3C, 0x24,
	0x01, 0x55, 0x1E, 0x3E, 0x36, 0x3B, 0x33, 0x41, 0x39, 0x21, 0x1F, 0x35,
	0x59, 0x13, 0x16, 0x1E, 0x31, 0x02, 0x06, 0x0D, 0x59, 0x31, 0x27, 0x2E,
	0x2D, 0x08, 0x04, 0x5C, 0x09, 0x32, 0x34, 0x05, 0x3E, 0x20, 0x23, 0x28,
	0x00, 0x28, 0x2A, 0x36, 0x22, 0x04, 0x03, 0x20, 0x2E, 0x0B, 0x38, 0x23,
	0x1C, 0x2F, 0x0A, 0x32, 0x39, 0x3E, 0x30, 0x15, 0x23, 0x3C, 0x28, 0x03,
	0x3A, 0x19, 0x3B, 0x05, 0x2F, 0x59, 0x4E, 0x21, 0x2D, 0x15, 0x36, 0x18,
	0x5A, 0x3F, 0x05, 0x47, 0x2A, 0x09, 0x2A, 0x36, 0x3D, 0x55, 0x24, 0x32,
	0x14, 0x07, 0x19, 0x16, 0x2A, 0x12, 0x3A, 0x59, 0x09, 0x27, 0x18, 0x2B,
	0x3B, 0x19, 0x13, 0x23, 0x05, 0x14, 0x2B, 0x5D, 0x20, 0x54, 0x05, 0x0D,
	0x00, 0x26, 0x0B, 0x0A, 0x34, 0x3B, 0x73, 0x0F, 0x27, 0x3C, 0x5F, 0x21,
	0x0F, 0x2C, 0x0C, 0x58, 0x03, 0x29, 0x34, 0x0D, 0x0D, 0x30, 0x0E, 0x51,
	0x2B, 0x0F, 0x7A, 0x29, 0x27, 0x2D, 0x3B, 0x3A, 0x04, 0x16, 0x36, 0x3B,
	0x21, 0x47, 0x08, 0x2D, 0x13, 0x71, 0x3D, 0x29, 0x59, 0x25, 0x69, 0x5D,
	0x57, 0x5F, 0x0A, 0x36, 0x14, 0x30, 0x5B, 0x0F, 0x33, 0x18, 0x39, 0x1E,
	0x09, 0x1A, 0x54, 0x29, 0x1F, 0x2E, 0x11, 0x55, 0x09, 0x21, 0x19, 0x2A,
	0x0D, 0x29, 0x3D, 0x29, 0x05, 0x5F, 0x39, 0x45, 0x09, 0x2F, 0x20, 0x2A,
	0x3D, 0x18, 0x2A, 0x1E, 0x2C, 0x34, 0x12, 0x75, 0x3F, 0x2A, 0x04, 0x3E,
	0x34, 0x3A, 0x25, 0x24, 0x01, 0x0B, 0x38, 0x03, 0x03, 0x40, 0x00, 0x2E,
	0x33, 0x00, 0x39, 0x76, 0x1F, 0x11, 0x17, 0x0A, 0x34, 0x36, 0x17, 0x37,
	0x00, 0x35, 0x38, 0x17, 0x21, 0x40, 0x2F, 0x55, 0x24, 0x5C, 0x5E, 0x24,
	0x54, 0x0B, 0x0A, 0x3B, 0x2A, 0x1A, 0x59, 0x07, 0x5F, 0x20, 0x55, 0x12,
	0x0A, 0x2E, 0x21, 0x27, 0x52, 0x20, 0x08, 0x06, 0x22, 0x51, 0x1C, 0x29,
	0x37, 0x3E, 0x52, 0x56, 0x5C, 0x03, 0x1C, 0x06, 0x23, 0x18, 0x08, 0x1C,
	0x4A, 0x06, 0x06, 0x25, 0x36, 0x0A, 0x38, 0x28, 0x27, 0x16, 0x2E, 0x09,
	0x23, 0x0D, 0x07, 0x2F, 0x24, 0x2A, 0x3B, 0x5D, 0x13, 0x3B, 0x2C, 0x0D,
	0x3E, 0x50, 0x5D, 0x0C, 0x1B, 0x5B, 0x09, 0x06, 0x00, 0x38, 0x06, 0x12,
	0x21, 0x26, 0x72, 0x09, 0x16, 0x17, 0x04, 0x14, 0x58, 0x51, 0x3B, 0x23,
	0x34, 0x08, 0x20, 0x36, 0x29, 0x21, 0x25, 0x34, 0x1E, 0x19, 0x6D, 0x58,
	0x15, 0x22, 0x44, 0x75, 0x01, 0x00, 0x2D, 0x00, 0x26, 0x5C, 0x23, 0x05,
	0x5B, 0x17, 0x20, 0x2E, 0x23, 0x26, 0x17, 0x5F, 0x0E, 0x3D, 0x5B, 0x11,
	0x09, 0x29, 0x2B, 0x04, 0x2B, 0x27, 0x03, 0x20, 0x03, 0x26, 0x22, 0x0A,
	0x56, 0x3D, 0x34, 0x5D, 0x2B, 0x1A, 0x04, 0x31, 0x09, 0x2C, 0x45, 0x58,
	0x73, 0x3D, 0x02, 0x3F, 0x20, 0x13, 0x1B, 0x11, 0x26, 0x5F, 0x15, 0x19,
	0x3B, 0x1B, 0x5A, 0x0C, 0x3E, 0x05, 0x25, 0x11, 0x75, 0x27, 0x55, 0x3F,
	0x09, 0x29, 0x3A, 0x16, 0x06, 0x19, 0x08, 0x2A, 0x14, 0x1D, 0x32, 0x27,
	0x18, 0x35, 0x04, 0x02, 0x20, 0x24, 0x06, 0x18, 0x1A, 0x38, 0x04, 0x30,
	0x2D, 0x58, 0x17, 0x2F, 0x26, 0x1B, 0x0C, 0x07, 0x35, 0x26, 0x37, 0x2D,
	0x01, 0x47, 0x54, 0x05, 0x23, 0x1B, 0x1F, 0x38, 0x41, 0x53, 0x33, 0x5D,
	0x35, 0x36, 0x0A, 0x13, 0x19, 0x06, 0x3A, 0x22, 0x74, 0x5E, 0x4A, 0x3B,
	0x40, 0x35, 0x08, 0x38, 0x19, 0x2D, 0x0A, 0x00, 0x1B, 0x1C, 0x09, 0x2E,
	0x43, 0x04, 0x5E, 0x21, 0x7A, 0x5F, 0x29, 0x01, 0x09, 0x2D, 0x20, 0x36,
	0x3A, 0x0F, 0x01, 0x2D, 0x39, 0x27, 0x2D, 0x77, 0x5E, 0x09, 0x2B, 0x52,
	0x17, 0x1F, 0x58, 0x25, 0x39, 0x31, 0x22, 0x54, 0x45, 0x3A, 0x77, 0x16,
	0x55, 0x01, 0x29, 0x0F, 0x1C, 0x0B, 0x03, 0x5D, 0x0B, 0x3E, 0x51, 0x0A,
	0x08, 0x25, 0x2F, 0x4E, 0x2A, 0x5B, 0x3A, 0x03, 0x38, 0x23, 0x5E, 0x75,
	0x2A, 0x1B, 0x3C, 0x31, 0x2B, 0x15, 0x2E, 0x04, 0x5A, 0x05, 0x02, 0x24,
	0x38, 0x39, 0x21, 0x3F, 0x00, 0x07, 0x31, 0x31, 0x2F, 0x0B, 0x07, 0x0F,
	0x25, 0x38, 0x2F, 0x03, 0x3D, 0x1A, 0x26, 0x0B, 0x5C, 0x03, 0x2B, 0x3D,
	0x14, 0x1A, 0x08, 0x37, 0x1B, 0x11, 0x56, 0x23, 0x07, 0x03, 0x39, 0x1B,
	0x21, 0x29, 0x16, 0x2D, 0x37, 0x31, 0x73, 0x21, 0x18, 0x58, 0x2D, 0x3B,
	0x1D, 0x27, 0x57, 0x59, 0x1B, 0x1C, 0x52, 0x1D, 0x25, 0x73, 0x25, 0x31,
	0x09, 0x31, 0x24, 0x29, 0x2A, 0x5E, 0x07, 0x20, 0x2F, 0x00, 0x3C, 0x13,
	0x35, 0x24, 0x2A, 0x1F, 0x07, 0x07, 0x14, 0x34, 0x3C, 0x12, 0x10, 0x0D,
	0x15, 0x09, 0x1D, 0x2E, 0x18, 0x0E, 0x08, 0x26, 0x06, 0x3E, 0x10, 0x57,
	0x1A, 0x2B, 0x26, 0x07, 0x09, 0x21, 0x08, 0x3E, 0x10, 0x09, 0x0F, 0x05,
	0x05, 0x4E, 0x41, 0x1A, 0x37, 0x2B, 0x53, 0x1C, 0x18, 0x11, 0x3E, 0x20,
	0x28, 0x5B, 0x74, 0x1D, 0x55, 0x3D, 0x3D, 0x04, 0x16, 0x2B, 0x22, 0x11,
	0x2E, 0x07, 0x29, 0x3F, 0x38, 0x06, 0x09, 0x51, 0x17, 0x02, 0x31, 0x1C,
	0x34, 0x07, 0x1E, 0x16, 0x2F, 0x33, 0x45, 0x13, 0x08, 0x2D, 0x2E, 0x22,
	0x5C, 0x31, 0x2A, 0x37, 0x5A, 0x5A, 0x34, 0x1B, 0x26, 0x2D, 0x58, 0x13,
	0x5D, 0x54, 0x02, 0x5F, 0x2F, 0x5F, 0x15, 0x3A, 0x5B, 0x15, 0x0B, 0x55,
	0x2B, 0x2A, 0x05, 0x0F, 0x27, 0x27, 0x0E, 0x28, 0x58, 0x05, 0x08, 0x0D,
	0x32, 0x28, 0x2F, 0x01, 0x5B, 0x7A, 0x0E, 0x29, 0x0A, 0x1F, 0x0B, 0x27,
	0x29, 0x0C, 0x07, 0x30, 0x03, 0x16, 0x0D, 0x19, 0x01, 0x38, 0x28, 0x1B,
	0x40, 0x05, 0x09, 0x29, 0x20, 0x06, 0x76, 0x0F, 0x15, 0x5E, 0x3D, 0x0C,
	0x28, 0x22, 0x5D, 0x29, 0x31, 0x0F, 0x1B, 0x0A, 0x1C, 0x0B, 0x16, 0x20,
	0x29, 0x5B, 0x35, 0x22, 0x0C, 0x27, 0x38, 0x0C, 0x3B, 0x31, 0x0B, 0x11,
	0x35, 0x05, 0x16, 0x5A, 0x2C, 0x27, 0x54, 0x29, 0x5D, 0x5C, 0x05, 0x28,
	0x11, 0x1A, 0x44, 0x7B, 0x0B, 0x53, 0x07, 0x5C, 0x74, 0x59, 0x0F, 0x02,
	0x3C, 0x30, 0x1E, 0x0E, 0x26, 0x19, 0x38, 0x24, 0x2A, 0x27, 0x0D, 0x08,
	0x25, 0x20, 0x0B, 0x53, 0x35, 0x22, 0x18, 0x41, 0x31, 0x1B, 0x3F, 0x2C,
	0x18, 0x27, 0x6D, 0x1E, 0x0F, 0x08, 0x3F, 0x73, 0x3B, 0x25, 0x2D, 0x26,
	0x27, 0x1F, 0x08, 0x27, 0x02, 0x3A, 0x2E, 0x23, 0x5B, 0x58, 0x29, 0x1C,
	0x2D, 0x0A, 0x01, 0x14, 0x5F, 0x0E, 0x00, 0x27, 0x26, 0x34, 0x54, 0x5E,
	0x1D, 0x2A, 0x01, 0x2F, 0x2F, 0x0F, 0x15, 0x3D, 0x20, 0x24, 0x02, 0x23,
	0x27, 0x20, 0x0A, 0x0E, 0x1A, 0x22, 0x25, 0x57, 0x5F, 0x30, 0x24, 0x09,
	0x38, 0x26, 0x09, 0x0F, 0x10, 0x16, 0x1E, 0x7A, 0x3B, 0x58, 0x03, 0x0D,
	0x34, 0x24, 0x14, 0x1D, 0x2F, 0x72, 0x3F, 0x2C, 0x3D, 0x3D, 0x11, 0x01,
	0x55, 0x41, 0x1A, 0x3A, 0x2A, 0x09, 0x18, 0x12, 0x69, 0x06, 0x24, 0x5A,
	0x29, 0x24, 0x1E, 0x0D, 0x36, 0x33, 0x33, 0x5D, 0x28, 0x2B, 0x3E, 0x0E,
	0x5F, 0x2D, 0x00, 0x53, 0x70, 0x43, 0x0C, 0x22, 0x2C, 0x77, 0x23, 0x51,
	0x18, 0x0C, 0x25, 0x18, 0x33, 0x37, 0x03, 0x34, 0x47, 0x28, 0x1A, 0x19,
	0x6D, 0x0F, 0x36, 0x36, 0x5F, 0x0F, 0x39, 0x50, 0x28, 0x38, 0x17, 0x39,
	0x55, 0x1A, 0x25, 0x2C, 0x29, 0x05, 0x17, 0x11, 0x26, 0x5C, 0x06, 0x3E,
	0x1F, 0x34, 0x3D, 0x1B, 0x56, 0x09, 0x1A, 0x38, 0x2D, 0x34, 0x38, 0x11,
	0x3E, 0x57, 0x0C, 0x33, 0x32, 0x3F, 0x39, 0x20, 0x2D, 0x0E, 0x3F, 0x11,
	0x1E, 0x08, 0x20, 0x24, 0x4E, 0x3D, 0x13, 0x36, 0x16, 0x08, 0x5C, 0x26,
	0x0C, 0x24, 0x33, 0x41, 0x59, 0x37, 0x0F, 0x24, 0x3A, 0x3A, 0x2E, 0x5B,
	0x54, 0x26, 0x26, 0x0F, 0x1C, 0x08, 0x0C, 0x59, 0x71, 0x59, 0x33, 0x3E,
	0x1C, 0x29, 0x1A, 0x00, 0x09, 0x28, 0x76, 0x34, 0x20, 0x39, 0x04, 0x08,
	0x2E, 0x0D, 0x09, 0x3C, 0x04, 0x35, 0x04, 0x5E, 0x20, 0x0B, 0x34, 0x52,
	0x07, 0x0C, 0x16, 0x3D, 0x25, 0x06, 0x3D, 0x13, 0x00, 0x00, 0x2D, 0x5E,
	0x69, 0x2A, 0x28, 0x29, 0x53, 0x26, 0x3F, 0x07, 0x3D, 0x1A, 0x2E, 0x47,
	0x03, 0x28, 0x11, 0x7B, 0x3F, 0x2F, 0x0B, 0x05, 0x69, 0x03, 0x36, 0x0F,
	0x0E, 0x30, 0x5D, 0x57, 0x00, 0x09, 0x7B, 0x5A, 0x26, 0x59, 0x24, 0x7A,
	0x1F, 0x0B, 0x09, 0x58, 0x76, 0x3B, 0x53, 0x3F, 0x40, 0x72, 0x5E, 0x23,
	0x26, 0x0D, 0x0C, 0x03, 0x12, 0x3D, 0x28, 0x00, 0x04, 0x11, 0x37, 0x2A,
	0x7A, 0x2E, 0x13, 0x03, 0x1F, 0x05, 0x47, 0x57, 0x1B, 0x03, 0x2B, 0x3B,
	0x51, 0x5A, 0x1F, 0x77, 0x22, 0x29, 0x1A, 0x08, 0x77, 0x5D, 0x06, 0x14,
	0x28, 0x28, 0x16, 0x50, 0x38, 0x04, 0x0F, 0x39, 0x19, 0x03, 0x04, 0x2E,
	0x3D, 0x10, 0x57, 0x00, 0x37, 0x22, 0x59, 0x01, 0x18, 0x25, 0x1B, 0x26,
	0x3D, 0x1B, 0x33, 0x58, 0x18, 0x3C, 0x0F, 0x26, 0x5A, 0x07, 0x1B, 0x1D,
	0x37, 0x19, 0x20, 0x5F, 0x22, 0x03, 0x5E, 0x15, 0x26, 0x21, 0x76, 0x14,
	0x58, 0x59, 0x0E, 0x74, 0x2E, 0x27, 0x00, 0x25, 0x2F, 0x58, 0x2B, 0x5F,
	0x19, 0x03, 0x3C, 0x32, 0x17, 0x1F, 0x18, 0x2E, 0x13, 0x0A, 0x58, 0x69,
	0x24, 0x56, 0x07, 0x22, 0x1B, 0x26, 0x17, 0x3D, 0x08, 0x14, 0x5B, 0x0B,
	0x3E, 0x3C, 0x03, 0x29, 0x00, 0x21, 0x58, 0x00, 0x09, 0x50, 0x0F, 0x29,
	0x37, 0x0D, 0x51, 0x5E, 0x3F, 0x25, 0x5D, 0x04, 0x02, 0x33, 0x09, 0x43,
	0x55, 0x2F, 0x3E, 0x06, 0x1F, 0x2A, 0x57, 0x06, 0x29, 0x38, 0x0E, 0x17,
	0x07, 0x76, 0x0E, 0x12, 0x1E, 0x1D, 0x73, 0x1E, 0x35, 0x34, 0x20, 0x21,
	0x2E, 0x58, 0x38, 0x3E, 0x0C, 0x5A, 0x14, 0x1E, 0x5A, 0x35, 0x24, 0x50,
	0x5F, 0x09, 0x2D, 0x35, 0x03, 0x00, 0x09, 0x35, 0x04, 0x31, 0x5C, 0x23,
	0x13, 0x0A, 0x2E, 0x59, 0x5B, 0x2A, 0x27, 0x24, 0x57, 0x1E, 0x0F, 0x0A,
	0x2D, 0x34, 0x5F, 0x23, 0x38, 0x58, 0x0F, 0x1F, 0x2C, 0x19, 0x0A, 0x1E,
	0x00, 0x38, 0x5F, 0x24, 0x0F, 0x2F, 0x0F, 0x1F, 0x2E, 0x1D, 0x5E, 0x3A,
	0x21, 0x59, 0x3A, 0x1D, 0x72, 0x27, 0x3B, 0x3E, 0x24, 0x16, 0x5B, 0x37,
	0x04, 0x58, 0x15, 0x1E, 0x29, 0x58, 0x05, 0x77, 0x1D, 0x52, 0x57, 0x3F,
	0x34, 0x15, 0x06, 0x29, 0x23, 0x04, 0x1B, 0x3B, 0x28, 0x06, 0x17, 0x1D,
	0x20, 0x17, 0x38, 0x77, 0x2F, 0x08, 0x0A, 0x29, 0x0F, 0x55, 0x25, 0x58,
	0x28, 0x3B, 0x2D, 0x0F, 0x2B, 0x53, 0x1A, 0x2E, 0x51, 0x59, 0x06, 0x72,
	0x2B, 0x34, 0x45, 0x22, 0x37, 0x23, 0x18, 0x2D, 0x1D, 0x28, 0x28, 0x14,
	0x2A, 0x32, 0x33, 0x5B, 0x32, 0x1D, 0x3A, 0x2E, 0x2E, 0x2E, 0x1C, 0x28,
	0x06, 0x09, 0x55, 0x5E, 0x59, 0x2D, 0x15, 0x35, 0x5B, 0x22, 0x36, 0x38,
	0x51, 0x27, 0x1F, 0x2F, 0x27, 0x2D, 0x21, 0x5A, 0x18, 0x2E, 0x16, 0x2A,
	0x1D, 0x15, 0x0B, 0x24, 0x5C, 0x3C, 0x16, 0x2B, 0x29, 0x2A, 0x21, 0x37,
	0x0D, 0x09, 0x57, 0x3E, 0x25, 0x2D, 0x12, 0x21, 0x5F, 0x34, 0x20, 0x28,
	0x1B, 0x26, 0x06, 0x09, 0x2A, 0x25, 0x5D, 0x15, 0x2F, 0x14, 0x25, 0x38,
	0x3B, 0x3D, 0x2D, 0x29, 0x2C, 0x33, 0x29, 0x55, 0x02, 0x2D, 0x7A, 0x35,
	0x0C, 0x3D, 0x5F, 0x17, 0x14, 0x05, 0x03, 0x40, 0x14, 0x0B, 0x2B, 0x16,
	0x1C, 0x7A, 0x01, 0x55, 0x0D, 0x09, 0x2D, 0x03, 0x29, 0x38, 0x1C, 0x12,
	0x02, 0x30, 0x28, 0x3B, 0x0A, 0x16, 0x2E, 0x1A, 0x1A, 0x74, 0x1E, 0x04,
	0x2F, 0x2D, 0x32, 0x2E, 0x19, 0x37, 0x5B, 0x70, 0x1F, 0x16, 0x5E, 0x1A,
	0x31, 0x5F, 0x10, 0x2B, 0x33, 0x10, 0x04, 0x2B, 0x09, 0x20, 0x05, 0x43,
	0x09, 0x29, 0x1D, 0x31, 0x06, 0x1B, 0x08, 0x5C, 0x37, 0x5C, 0x15, 0x1E,
	0x2D, 0x1B, 0x07, 0x55, 0x0D, 0x0D, 0x2E, 0x24, 0x23, 0x0C, 0x3A, 0x72,
	0x05, 0x2E, 0x16, 0x5A, 0x76, 0x3C, 0x4A, 0x2F, 0x29, 0x73, 0x3C, 0x03,
	0x03, 0x2E, 0x29, 0x5A, 0x16, 0x3B, 0x06, 0x24, 0x3D, 0x25, 0x0B, 0x44,
	0x0B, 0x06, 0x52, 0x17, 0x19, 0x20, 0x5E, 0x35, 0x34, 0x3A, 0x14, 0x0D,
	0x00, 0x3A, 0x33, 0x7A, 0x1D, 0x2F, 0x41, 0x21, 0x37, 0x1F, 0x2A, 0x5E,
	0x22, 0x26, 0x5E, 0x15, 0x25, 0x44, 0x2B, 0x20, 0x14, 0x0A, 0x28, 0x7A,
	0x2D, 0x11, 0x04, 0x33, 0x2D, 0x55, 0x0A, 0x1A, 0x26, 0x30, 0x29, 0x30,
	0x00, 0x23, 0x11, 0x5E, 0x0C, 0x5A, 0x06, 0x04, 0x03, 0x22, 0x28, 0x1C,
	0x03, 0x38, 0x29, 0x28, 0x18, 0x0D, 0x3D, 0x55, 0x37, 0x02, 0x05, 0x0F,
	0x37, 0x1A, 0x32, 0x05, 0x5D, 0x39, 0x29, 0x28, 0x25, 0x0E, 0x13, 0x17,
	0x01, 0x76, 0x26, 0x58, 0x45, 0x1A, 0x30, 0x25, 0x3B, 0x21, 0x5C, 0x71,
	0x3E, 0x32, 0x5E, 0x1F, 0x24, 0x59, 0x31, 0x00, 0x2D, 0x3A, 0x2E, 0x22,
	0x5E, 0x2D, 0x7A, 0x2E, 0x2F, 0x5E, 0x2E, 0x2A, 0x21, 0x50, 0x3A, 0x5C,
	0x76, 0x28, 0x51, 0x39, 0x2A, 0x1B, 0x0D, 0x32, 0x2D, 0x08, 0x18, 0x58,
	0x31, 0x0A, 0x11, 0x03, 0x2D, 0x03, 0x56, 0x3B, 0x13, 0x02, 0x00, 0x28,
	0x0E, 0x04, 0x0F, 0x10, 0x59, 0x2E, 0x1B, 0x1B, 0x0A, 0x59, 0x5F, 0x06,
	0x0A, 0x2A, 0x5B, 0x20, 0x75, 0x5F, 0x56, 0x1A, 0x3C, 0x28, 0x1A, 0x2F,
	0x0C, 0x19, 0x1A, 0x0E, 0x2C, 0x3E, 0x01, 0x1A, 0x18, 0x08, 0x20, 0x04,
	0x32, 0x3D, 0x3B, 0x41, 0x1A, 0x2E, 0x16, 0x0C, 0x37, 0x20, 0x08, 0x15,
	0x2D, 0x0B, 0x09, 0x0B, 0x2A, 0x25, 0x5F, 0x5E, 0x28, 0x38, 0x13, 0x0D,
	0x01, 0x2D, 0x08, 0x16, 0x38, 0x22, 0x23, 0x05, 0x56, 0x00, 0x2C, 0x75,
	0x24, 0x27, 0x26, 0x3A, 0x0A, 0x2E, 0x25, 0x3A, 0x2A, 0x3A, 0x05, 0x23,
	0x1F, 0x31, 0x15, 0x3F, 0x38, 0x06, 0x44, 0x35, 0x1A, 0x4E, 0x2F, 0x0F,
	0x72, 0x0B, 0x52, 0x08, 0x07, 0x7B, 0x5F, 0x16, 0x41, 0x3C, 0x06, 0x5D,
	0x26, 0x5D, 0x11, 0x0E, 0x58, 0x28, 0x29, 0x26, 0x73, 0x0B, 0x32, 0x28,
	0x33, 0x17, 0x3F, 0x27, 0x26, 0x3A, 0x34, 0x35, 0x36, 0x1D, 0x38, 0x26,
	0x1F, 0x32, 0x0D, 0x3E, 0x2D, 0x1A, 0x06, 0x3A, 0x05, 0x07, 0x05, 0x50,
	0x01, 0x32, 0x2E, 0x39, 0x2F, 0x5D, 0x18, 0x1A, 0x14, 0x25, 0x37, 0x28,
	0x14, 0x2D, 0x0D, 0x5A, 0x22, 0x09, 0x0E, 0x0D, 0x39, 0x5C, 0x37, 0x05,
	0x07, 0x1F, 0x22, 0x15, 0x05, 0x22, 0x3C, 0x1B, 0x71, 0x3D, 0x28, 0x07,
	0x20, 0x3A, 0x0A, 0x00, 0x23, 0x59, 0x1A, 0x18, 0x59, 0x1A, 0x18, 0x2B,
	0x01, 0x34, 0x05, 0x59, 0x32, 0x22, 0x20, 0x03, 0x01, 0x14, 0x1A, 0x20,
	0x5C, 0x38, 0x14, 0x2D, 0x4E, 0x24, 0x11, 0x17, 0x1B, 0x55, 0x01, 0x3E,
	0x73, 0x5B, 0x36, 0x2F, 0x06, 0x2E, 0x2E, 0x22, 0x09, 0x5B, 0x28, 0x58,
	0x20, 0x2B, 0x05, 0x33, 0x1A, 0x0D, 0x34, 0x1C, 0x1A, 0x5D, 0x14, 0x36,
	0x1E, 0x70, 0x43, 0x09, 0x00, 0x27, 0x06, 0x2A, 0x12, 0x38, 0x5A, 0x2A,
	0x5F, 0x16, 0x19, 0x38, 0x2D, 0x43, 0x20, 0x59, 0x59, 0x28, 0x2E, 0x2B,
	0x1D, 0x1F, 0x0C, 0x3B, 0x24, 0x2B, 0x20, 0x20, 0x58, 0x30, 0x2F, 0x05,
	0x26, 0x16, 0x2A, 0x58, 0x08, 0x17, 0x3B, 0x2E, 0x5F, 0x1F, 0x36, 0x5E,
	0x14, 0x2C, 0x53, 0x09, 0x2B, 0x15, 0x5D, 0x0C, 0x05, 0x1E, 0x2A, 0x3D,
	0x33, 0x0B, 0x27, 0x06, 0x07, 0x3C, 0x6D, 0x3F, 0x57, 0x2F, 0x31, 0x0E,
	0x0E, 0x0F, 0x3A, 0x01, 0x34, 0x24, 0x32, 0x57, 0x1B, 0x26, 0x16, 0x0E,
	0x16, 0x06, 0x31, 0x2F, 0x2C, 0x3C, 0x0C, 0x20, 0x3A, 0x2C, 0x58, 0x12,
	0x3A, 0x1D, 0x30, 0x14, 0x27, 0x27, 0x2B, 0x50, 0x04, 0x2C, 0x13, 0x28,
	0x15, 0x14, 0x13, 0x07, 0x15, 0x17, 0x56, 0x1D, 0x01, 0x38, 0x20, 0x2A,
	0x01, 0x20, 0x59, 0x27, 0x17, 0x27, 0x3B, 0x24, 0x0F, 0x2F, 0x22, 0x3B,
	0x23, 0x30, 0x39, 0x40, 0x3B, 0x3F, 0x0F, 0x09, 0x39, 0x32, 0x3D, 0x24,
	0x36, 0x19, 0x3A, 0x3C, 0x0D, 0x2B, 0x39, 0x15, 0x5F, 0x51, 0x16, 0x1A,
	0x01, 0x0B, 0x17, 0x0F, 0x40, 0x23, 0x43, 0x0C, 0x3F, 0x3B, 0x31, 0x39,
	0x2E, 0x17, 0x03, 0x11, 0x28, 0x19, 0x18, 0x1F, 0x15, 0x18, 0x07, 0x14,
	0x5E, 0x15, 0x06, 0x53, 0x2D, 0x1E, 0x6D, 0x18, 0x22, 0x06, 0x22, 0x06,
	0x01, 0x32, 0x5E, 0x26, 0x7A, 0x5F, 0x27, 0x18, 0x20, 0x2A, 0x06, 0x0D,
	0x37, 0x52, 0x17, 0x39, 0x0D, 0x2F, 0x3A, 0x72, 0x20, 0x32, 0x5E, 0x07,
	0x3B, 0x2B, 0x53, 0x36, 0x32, 0x06, 0x08, 0x2D, 0x1B, 0x00, 0x75, 0x25,
	0x36, 0x58, 0x28, 0x07, 0x5A, 0x33, 0x22, 0x5C, 0x0B, 0x1F, 0x31, 0x19,
	0x22, 0x12, 0x0F, 0x26, 0x37, 0x3F, 0x38, 0x0F, 0x24, 0x5E, 0x08, 0x75,
	0x36, 0x28, 0x07, 0x5C, 0x05, 0x09, 0x2D, 0x2D, 0x07, 0x72, 0x2E, 0x31,
	0x04, 0x22, 0x0E, 0x0A, 0x15, 0x1B, 0x2A, 0x2C, 0x23, 0x3B, 0x45, 0x38,
	0x0C, 0x1C, 0x0C, 0x01, 0x23, 0x37, 0x0B, 0x58, 0x36, 0x58, 0x21, 0x3D,
	0x22, 0x1C, 0x22, 0x12, 0x3C, 0x24, 0x01, 0x0C, 0x01, 0x38, 0x31, 0x5C,
	0x0C, 0x1B, 0x0F, 0x28, 0x19, 0x23, 0x13, 0x3B, 0x57, 0x2B, 0x3F, 0x27,
	0x19, 0x0B, 0x59, 0x05, 0x09, 0x39, 0x11, 0x2C, 0x5F, 0x25, 0x04, 0x57,
	0x05, 0x25, 0x25, 0x3C, 0x24, 0x22, 0x3E, 0x08, 0x3C, 0x0D, 0x20, 0x2F,
	0x17, 0x5A, 0x38, 0x14, 0x02, 0x34, 0x19, 0x56, 0x5D, 0x26, 0x69, 0x25,
	0x15, 0x01, 0x25, 0x31, 0x55, 0x14, 0x5C, 0x2A, 0x2F, 0x1D, 0x20, 0x5B,
	0x29, 0x2F, 0x55, 0x07, 0x1D, 0x2A, 0x11, 0x1A, 0x10, 0x19, 0x2E, 0x1A,
	0x1C, 0x06, 0x18, 0x0E, 0x25, 0x3F, 0x02, 0x02, 0x32, 0x09, 0x2F, 0x31,
	0x21, 0x3F, 0x35, 0x03, 0x38, 0x37, 0x1C, 0x0D, 0x3F, 0x12, 0x2C, 0x01,
	0x1A, 0x26, 0x0F, 0x03, 0x0F, 0x08, 0x2E, 0x05, 0x0C, 0x13, 0x7B, 0x58,
	0x35, 0x1D, 0x22, 0x0A, 0x24, 0x11, 0x3F, 0x0C, 0x7A, 0x19, 0x53, 0x23,
	0x23, 0x74, 0x5C, 0x2C, 0x29, 0x1E, 0x77, 0x03, 0x08, 0x0B, 0x00, 0x1B,
	0x28, 0x56, 0x1C, 0x1D, 0x7B, 0x1B, 0x02, 0x3A, 0x01, 0x05, 0x3A, 0x03,
	0x5A, 0x26, 0x32, 0x02, 0x2E, 0x39, 0x2E, 0x2D, 0x47, 0x16, 0x01, 0x0A,
	0x71, 0x2E, 0x02, 0x04, 0x01, 0x23, 0x5A, 0x17, 0x59, 0x3F, 0x1B, 0x58,
	0x0E, 0x04, 0x3C, 0x25, 0x07, 0x3B, 0x1D, 0x07, 0x74, 0x3D, 0x52, 0x1E,
	0x26, 0x33, 0x1C, 0x02, 0x5C, 0x39, 0x36, 0x08, 0x10, 0x28, 0x26, 0x0D,
	0x14, 0x0A, 0x04, 0x21, 0x72, 0x3B, 0x3B, 0x5A, 0x2F, 0x2E, 0x07, 0x0C,
	0x5E, 0x02, 0x74, 0x1C, 0x19, 0x18, 0x58, 0x26, 0x20, 0x19, 0x3D, 0x2C,
	0x31, 0x59, 0x2A, 0x1F, 0x3C, 0x69, 0x47, 0x19, 0x24, 0x3B, 0x12, 0x04,
	0x06, 0x38, 0x5F, 0x24, 0x0B, 0x20, 0x3C, 0x19, 0x3B, 0x24, 0x19, 0x5A,
	0x1B, 0x28, 0x0A, 0x38, 0x58, 0x05, 0x32, 0x1B, 0x51, 0x1C, 0x33, 0x13,
	0x0F, 0x12, 0x3E, 0x1C, 0x2D, 0x23, 0x13, 0x26, 0x07, 0x03, 0x47, 0x4A,
	0x20, 0x2D, 0x74, 0x1C, 0x24, 0x37, 0x12, 0x2C, 0x5A, 0x3B, 0x38, 0x38,
	0x0B, 0x0A, 0x32, 0x38, 0x07, 0x00, 0x1E, 0x23, 0x1C, 0x26, 0x16, 0x38,
	0x55, 0x36, 0x40, 0x1B, 0x07, 0x1B, 0x0F, 0x13, 0x24, 0x0E, 0x27, 0x5F,
	0x27, 0x33, 0x23, 0x51, 0x3F, 0x0A, 0x28, 0x2E, 0x24, 0x18, 0x0D, 0x70,
	0x2A, 0x18, 0x23, 0x26, 0x15, 0x3E, 0x2A, 0x22, 0x19, 0x14, 0x1F, 0x09,
	0x1D, 0x2D, 0x75, 0x55, 0x0B, 0x37, 0x22, 0x04, 0x3F, 0x16, 0x1C, 0x26,
	0x73, 0x3A, 0x0B, 0x07, 0x5C, 0x3B, 0x15, 0x19, 0x22, 0x23, 0x2A, 0x35,
	0x06, 0x0C, 0x00, 0x37, 0x0E, 0x07, 0x01, 0x07, 0x09, 0x26, 0x35, 0x0D,
	0x23, 0x72, 0x20, 0x25, 0x02, 0x1E, 0x28, 0x2B, 0x0D, 0x2A, 0x5F, 0x38,
	0x0B, 0x2D, 0x5B, 0x3D, 0x2A, 0x18, 0x55, 0x1D, 0x3B, 0x35, 0x05, 0x2D,
	0x37, 0x1F, 0x2A, 0x28, 0x00, 0x19, 0x04, 0x14, 0x5C, 0x20, 0x09, 0x44,
	0x15, 0x1D, 0x04, 0x3B, 0x5D, 0x03, 0x3E, 0x2D, 0x3B, 0x1F, 0x11, 0x2F,
	0x52, 0x3C, 0x53, 0x08, 0x2F, 0x0D, 0x00, 0x07, 0x0D, 0x47, 0x17, 0x57,
	0x07, 0x09, 0x28, 0x33, 0x22, 0x05, 0x13, 0x0A, 0x53, 0x3F, 0x33, 0x03,
	0x2D, 0x56, 0x24, 0x3C, 0x01, 0x43, 0x0D, 0x5B, 0x2F, 0x70, 0x39, 0x2F,
	0x5B, 0x01, 0x14, 0x1C, 0x0A, 0x3E, 0x0C, 0x72, 0x3C, 0x27, 0x23, 0x33,
	0x75, 0x28, 0x56, 0x26, 0x18, 0x31, 0x07, 0x31, 0x04, 0x00, 0x06, 0x29,
	0x09, 0x1B, 0x04, 0x23, 0x09, 0x20, 0x22, 0x1F, 0x0A, 0x06, 0x13, 0x29,
	0x5A, 0x23, 0x16, 0x2C, 0x3B, 0x01, 0x3B, 0x0F, 0x22, 0x05, 0x58, 0x71,
	0x00, 0x07, 0x0D, 0x29, 0x3B, 0x04, 0x57, 0x28, 0x5E, 0x26, 0x59, 0x2C,
	0x25, 0x40, 0x0A, 0x2E, 0x25, 0x5C, 0x58, 0x37, 0x5D, 0x03, 0x3A, 0x1B,
	0x21, 0x20, 0x59, 0x3C, 0x38, 0x38, 0x25, 0x2A, 0x28, 0x18, 0x37, 0x1A,
	0x2B, 0x20, 0x28, 0x06, 0x08, 0x08, 0x3D, 0x28, 0x11, 0x1F, 0x55, 0x0C,
	0x40, 0x75, 0x06, 0x39, 0x5E, 0x1E, 0x23, 0x07, 0x28, 0x28, 0x18, 0x12,
	0x0A, 0x04, 0x21, 0x58, 0x35, 0x25, 0x2A, 0x00, 0x21, 0x09, 0x2E, 0x1B,
	0x36, 0x5E, 0x30, 0x3F, 0x03, 0x2A, 0x58, 0x01, 0x0D, 0x2A, 0x0D, 0x0A,
	0x37, 0x00, 0x05, 0x28, 0x29, 0x77, 0x02, 0x4A, 0x01, 0x01, 0x12, 0x08,
	0x17, 0x5A, 0x18, 0x27, 0x21, 0x59, 0x1A, 0x33, 0x13, 0x36, 0x12, 0x5E,
	0x11, 0x12, 0x25, 0x35, 0x58, 0x25, 0x18, 0x25, 0x00, 0x28, 0x23, 0x0F,
	0x43, 0x03, 0x1B, 0x2A, 0x03, 0x3B, 0x10, 0x2D, 0x2D, 0x0A, 0x05, 0x55,
	0x0C, 0x28, 0x0B, 0x01, 0x17, 0x23, 0x3B, 0x09, 0x58, 0x29, 0x0D, 0x0C,
	0x34, 0x0B, 0x0C, 0x37, 0x05, 0x35, 0x3F, 0x15, 0x2C, 0x5B, 0x30, 0x59,
	0x25, 0x17, 0x3D, 0x76, 0x22, 0x2F, 0x59, 0x01, 0x01, 0x1B, 0x36, 0x3A,
	0x21, 0x3A, 0x35, 0x03, 0x17, 0x58, 0x73, 0x3B, 0x25, 0x5B, 0x05, 0x13,
	0x14, 0x26, 0x3A, 0x5E, 0x09, 0x06, 0x2C, 0x07, 0x09, 0x6D, 0x1C, 0x4E,
	0x00, 0x44, 0x21, 0x43, 0x57, 0x5E, 0x2F, 0x27, 0x0D, 0x50, 0x26, 0x0E,
	0x06, 0x16, 0x56, 0x41, 0x26, 0x15, 0x55, 0x39, 0x27, 0x06, 0x6D, 0x1A,
	0x4E, 0x14, 0x5C, 0x34, 0x09, 0x35, 0x2C, 0x1D, 0x24, 0x59, 0x35, 0x5D,
	0x52, 0x06, 0x43, 0x0A, 0x22, 0x38, 0x2F, 0x28, 0x05, 0x56, 0x3F, 0x00,
	0x0E, 0x53, 0x07, 0x2A, 0x29, 0x01, 0x36, 0x0C, 0x2E, 0x11, 0x3A, 0x37,
	0x03, 0x0F, 0x12, 0x23, 0x28, 0x21, 0x1D, 0x0F, 0x26, 0x32, 0x57, 0x2A,
	0x11, 0x3D, 0x4E, 0x41, 0x3E, 0x72, 0x01, 0x25, 0x37, 0x2E, 0x2E, 0x5F,
	0x02, 0x28, 0x02, 0x11, 0x0F, 0x04, 0x0B, 0x38, 0x71, 0x2E, 0x30, 0x02,
	0x0D, 0x15, 0x09, 0x2A, 0x16, 0x5D, 0x28, 0x2E, 0x13, 0x56, 0x11, 0x33,
	0x39, 0x2F, 0x5C, 0x44, 0x37, 0x04, 0x04, 0x0A, 0x00, 0x0D, 0x15, 0x57,
	0x3C, 0x09, 0x71, 0x00, 0x16, 0x00, 0x38, 0x29, 0x54, 0x0A, 0x0B, 0x3C,
	0x24, 0x3C, 0x31, 0x21, 0x11, 0x11, 0x16, 0x54, 0x3C, 0x18, 0x29, 0x14,
	0x38, 0x25, 0x27, 0x77, 0x24, 0x07, 0x04, 0x1B, 0x2E, 0x1E, 0x19, 0x3B,
	0x39, 0x33, 0x08, 0x32, 0x5A, 0x40, 0x00, 0x2A, 0x00, 0x20, 0x3B, 0x2A,
	0x08, 0x57, 0x20, 0x0C, 0x7A, 0x3E, 0x04, 0x2D, 0x07, 0x17, 0x19, 0x02,
	0x5E, 0x39, 0x13, 0x35, 0x2A, 0x21, 0x53, 0x69, 0x3A, 0x36, 0x04, 0x39,
	0x15, 0x3C, 0x1B, 0x38, 0x29, 0x7A, 0x16, 0x33, 0x3D, 0x52, 0x30, 0x1F,
	0x09, 0x20, 0x28, 0x35, 0x3D, 0x33, 0x34, 0x2A, 0x13, 0x23, 0x10, 0x28,
	0x08, 0x01, 0x1A, 0x55, 0x3C, 0x2E, 0x04, 0x0E, 0x2E, 0x1E, 0x01, 0x00,
	0x09, 0x31, 0x1B, 0x5B, 0x03, 0x1A, 0x2C, 0x19, 0x0E, 0x03, 0x14, 0x35,
	0x1A, 0x20, 0x36, 0x3A, 0x2C, 0x1B, 0x5B, 0x20, 0x5B, 0x31, 0x25, 0x02,
	0x34, 0x47, 0x25, 0x0A, 0x27, 0x7B, 0x23, 0x4A, 0x19, 0x3F, 0x07, 0x2E,
	0x0C, 0x1B, 0x1A, 0x2E, 0x05, 0x0B, 0x0D, 0x39, 0x18, 0x5E, 0x15, 0x28,
	0x2E, 0x2A, 0x05, 0x11, 0x06, 0x22, 0x2E, 0x27, 0x0C, 0x2C, 0x22, 0x28,
	0x43, 0x51, 0x5D, 0x2E, 0x2A, 0x5C, 0x0D, 0x3F, 0x25, 0x13, 0x5C, 0x30,
	0x3E, 0x27, 0x21, 0x3E, 0x05, 0x07, 0x26, 0x0C, 0x2D, 0x38, 0x3B, 0x1B,
	0x2A, 0x1F, 0x29, 0x28, 0x26, 0x01, 0x06, 0x33, 0x2C, 0x1C, 0x0D, 0x19,
	0x10, 0x26, 0x0E, 0x0E, 0x28, 0x17, 0x1E, 0x1C, 0x30, 0x08, 0x06, 0x41,
	0x2D, 0x23, 0x5A, 0x26, 0x16, 0x06, 0x07, 0x58, 0x22, 0x39, 0x32, 0x0C,
	0x39, 0x19, 0x25, 0x52, 0x10, 0x04, 0x05, 0x2D, 0x0F, 0x06, 0x1B, 0x17,
	0x34, 0x40, 0x0E, 0x03, 0x29, 0x07, 0x01, 0x77, 0x47, 0x0A, 0x1E, 0x21,
	0x36, 0x3F, 0x10, 0x14, 0x1B, 0x0E, 0x01, 0x2F, 0x24, 0x09, 0x77, 0x27,
	0x2F, 0x2B, 0x22, 0x36, 0x1E, 0x04, 0x3F, 0x52, 0x6D, 0x2A, 0x16, 0x1A,
	0x20, 0x17, 0x0F, 0x34, 0x22, 0x39, 0x7A, 0x22, 0x26, 0x03, 0x22, 0x10,
	0x5C, 0x33, 0x2D, 0x27, 0x17, 0x29, 0x2C, 0x23, 0x2A, 0x08, 0x3A, 0x05,
	0x18, 0x32, 0x23, 0x35, 0x26, 0x02, 0x1B, 0x09, 0x3B, 0x33, 0x07, 0x18,
	0x7A, 0x09, 0x18, 0x3E, 0x18, 0x06, 0x3B, 0x28, 0x34, 0x23, 0x03, 0x20,
	0x28, 0x28, 0x3B, 0x31, 0x25, 0x30, 0x57, 0x0A, 0x25, 0x34, 0x0C, 0x5B,
	0x19, 0x73, 0x1E, 0x2D, 0x0F, 0x1D, 0x08, 0x5B, 0x37, 0x5F, 0x29, 0x77,
	0x1E, 0x26, 0x1E, 0x3A, 0x3B, 0x3A, 0x2F, 0x05, 0x31, 0x1B, 0x43, 0x0D,
	0x41, 0x04, 0x10, 0x3B, 0x34, 0x01, 0x2E, 0x09, 0x47, 0x50, 0x21, 0x19,
	0x70, 0x58, 0x31, 0x2D, 0x1B, 0x07, 0x55, 0x0D, 0x09, 0x3B, 0x32, 0x2B,
	0x4E, 0x3A, 0x44, 0x69, 0x0B, 0x13, 0x45, 0x28, 0x30, 0x23, 0x57, 0x16,
	0x13, 0x03, 0x00, 0x10, 0x3C, 0x27, 0x26, 0x18, 0x59, 0x3D, 0x0E, 0x13,
	0x04, 0x4E, 0x3E, 0x11, 0x31, 0x0B, 0x15, 0x28, 0x0C, 0x76, 0x28, 0x2C,
	0x37, 0x5E, 0x1B, 0x1A, 0x28, 0x05, 0x13, 0x1B, 0x16, 0x31, 0x03, 0x5C,
	0x01, 0x0F, 0x23, 0x39, 0x0F, 0x1A, 0x3E, 0x0C, 0x5F, 0x1D, 0x72, 0x0D,
	0x24, 0x29, 0x24, 0x03, 0x3C, 0x14, 0x45, 0x39, 0x08, 0x04, 0x0E, 0x2B,
	0x39, 0x04, 0x3E, 0x17, 0x19, 0x24, 0x31, 0x27, 0x2E, 0x3D, 0x3C, 0x21,
	0x2E, 0x12, 0x34, 0x02, 0x7A, 0x3D, 0x05, 0x5A, 0x01, 0x21, 0x39, 0x56,
	0x0F, 0x2F, 0x10, 0x3E, 0x4E, 0x25, 0x2C, 0x2E, 0x59, 0x32, 0x0B, 0x5B,
	0x12, 0x5A, 0x09, 0x37, 0x20, 0x6D, 0x22, 0x59, 0x1A, 0x13, 0x77, 0x05,
	0x51, 0x3F, 0x03, 0x71, 0x1E, 0x55, 0x01, 0x1D, 0x72, 0x35, 0x1B, 0x16,
	0x3B, 0x7B, 0x01, 0x10, 0x41, 0x3C, 0x6D, 0x18, 0x15, 0x5D, 0x0A, 0x3A,
	0x5A, 0x53, 0x16, 0x32, 0x06, 0x59, 0x37, 0x01, 0x0A, 0x0C, 0x18, 0x18,
	0x06, 0x01, 0x18, 0x0F, 0x33, 0x25, 0x2E, 0x26, 0x2B, 0x0C, 0x00, 0x02,
	0x7A, 0x5B, 0x0D, 0x0F, 0x06, 0x14, 0x36, 0x53, 0x26, 0x03, 0x05, 0x0B,
	0x08, 0x3D, 0x3E, 0x08, 0x18, 0x16, 0x1D, 0x38, 0x71, 0x5B, 0x36, 0x2F,
	0x0A, 0x1A, 0x14, 0x2A, 0x00, 0x1F, 0x01, 0x25, 0x16, 0x41, 0x1D, 0x09,
	0x28, 0x2F, 0x1E, 0x03, 0x35, 0x59, 0x24, 0x1D, 0x53, 0x17, 0x5E, 0x36,
	0x45, 0x05, 0x73, 0x0D, 0x36, 0x3F, 0x04, 0x37, 0x5F, 0x18, 0x36, 0x2A,
	0x30, 0x26, 0x3B, 0x1F, 0x29, 0x04, 0x5D, 0x4E, 0x2C, 0x2E, 0x21, 0x20,
	0x00, 0x21, 0x0A, 0x76, 0x02, 0x2A, 0x36, 0x00, 0x0A, 0x3F, 0x35, 0x2C,
	0x06, 0x15, 0x3A, 0x50, 0x09, 0x23, 0x69, 0x3E, 0x36, 0x3F, 0x5A, 0x2B,
	0x2E, 0x1B, 0x1D, 0x1B, 0x1A, 0x55, 0x39, 0x1C, 0x0C, 0x31, 0x3D, 0x55,
	0x3B, 0x1C, 0x08, 0x18, 0x58, 0x41, 0x02, 0x74, 0x58, 0x05, 0x2A, 0x5D,
	0x73, 0x14, 0x50, 0x03, 0x0E, 0x1B, 0x2D, 0x14, 0x17, 0x44, 0x72, 0x5C,
	0x07, 0x17, 0x29, 0x25, 0x5E, 0x09, 0x5C, 0x19, 0x0B, 0x3D, 0x38, 0x14,
	0x5B, 0x10, 0x27, 0x13, 0x06, 0x2F, 0x32, 0x06, 0x06, 0x57, 0x13, 0x72,
	0x39, 0x18, 0x19, 0x38, 0x0A, 0x16, 0x2F, 0x5E, 0x06, 0x74, 0x2A, 0x14,
	0x37, 0x2A, 0x3B, 0x1A, 0x37, 0x28, 0x39, 0x29, 0x34, 0x29, 0x16, 0x08,
	0x36, 0x3F, 0x55, 0x2D, 0x02, 0x34, 0x01, 0x18, 0x38, 0x1A, 0x3B, 0x38,
	0x4E, 0x3F, 0x23, 0x33, 0x1F, 0x0F, 0x39, 0x00, 0x70, 0x0D, 0x2A, 0x17,
	0x05, 0x17, 0x3F, 0x50, 0x3D, 0x1B, 0x32, 0x3A, 0x30, 0x0A, 0x1A, 0x2E,
	0x54, 0x2B, 0x23, 0x1A, 0x30, 0x36, 0x32, 0x20, 0x31, 0x37, 0x47, 0x52,
	0x1E, 0x0F, 0x27, 0x24, 0x15, 0x1D, 0x1F, 0x23, 0x25, 0x0B, 0x1B, 0x0F,
	0x18, 0x5A, 0x36, 0x17, 0x5A, 0x7A, 0x2A, 0x2E, 0x58, 0x2C, 0x69, 0x09,
	0x06, 0x2F, 0x5D, 0x2F, 0x5D, 0x59, 0x24, 0x2E, 0x06, 0x16, 0x32, 0x24,
	0x23, 0x27, 0x39, 0x2B, 0x18, 0x11, 0x00, 0x06, 0x02, 0x25, 0x1D, 0x38,
	0x58, 0x39, 0x05, 0x27, 0x73, 0x1E, 0x4E, 0x0F, 0x04, 0x6D, 0x1A, 0x54,
	0x45, 0x3C, 0x36, 0x08, 0x56, 0x2C, 0x00, 0x1B, 0x25, 0x11, 0x18, 0x29,
	0x36, 0x25, 0x55, 0x5C, 0x20, 0x01, 0x5D, 0x0E, 0x24, 0x13, 0x06, 0x5B,
	0x50, 0x18, 0x5E, 0x16, 0x5D, 0x0F, 0x27, 0x26, 0x24, 0x3D, 0x2F, 0x5B,
	0x39, 0x0B, 0x08, 0x36, 0x23, 0x5B, 0x24, 0x1D, 0x23, 0x01, 0x07, 0x34,
	0x2E, 0x50, 0x02, 0x0F, 0x1B, 0x20, 0x0F, 0x36, 0x5B, 0x17, 0x1C, 0x37,
	0x2B, 0x0D, 0x33, 0x34, 0x56, 0x2B, 0x40, 0x28, 0x26, 0x0C, 0x07, 0x31,
	0x25, 0x3D, 0x16, 0x16, 0x5A, 0x74, 0x22, 0x09, 0x2D, 0x3C, 0x7B, 0x3F,
	0x34, 0x25, 0x3F, 0x72, 0x29, 0x55, 0x17, 0x58, 0x37, 0x1F, 0x00, 0x5E,
	0x24, 0x29, 0x23, 0x53, 0x02, 0x09, 0x25, 0x23, 0x2F, 0x34, 0x3E, 0x17,
	0x5F, 0x37, 0x56, 0x24, 0x15, 0x1D, 0x18, 0x28, 0x29, 0x16, 0x34, 0x2D,
	0x24, 0x3C, 0x2A, 0x1C, 0x11, 0x5F, 0x11, 0x20, 0x0D, 0x18, 0x38, 0x08,
	0x34, 0x55, 0x24, 0x28, 0x2D, 0x09, 0x01, 0x24, 0x3C, 0x01, 0x07, 0x5B,
	0x4E, 0x39, 0x3A, 0x15, 0x05, 0x58, 0x57, 0x38, 0x31, 0x29, 0x13, 0x28,
	0x0E, 0x2A, 0x15, 0x51, 0x02, 0x1C, 0x29, 0x22, 0x1B, 0x1C, 0x3F, 0x01,
	0x0B, 0x4E, 0x1A, 0x06, 0x34, 0x1E, 0x20, 0x1F, 0x06, 0x03, 0x14, 0x10,
	0x3D, 0x3A, 0x23, 0x47, 0x10, 0x23, 0x24, 0x00, 0x1F, 0x38, 0x1B, 0x1A,
	0x2A, 0x1D, 0x2A, 0x1E, 0x24, 0x12, 0x29, 0x34, 0x26, 0x02, 0x09, 0x47,
	0x39, 0x09, 0x05, 0x04, 0x26, 0x0F, 0x5D, 0x53, 0x05, 0x0A, 0x2B, 0x5F,
	0x1E, 0x0F, 0x38, 0x0E, 0x1D, 0x29, 0x76, 0x55, 0x27, 0x04, 0x25, 0x69,
	0x00, 0x23, 0x3A, 0x40, 0x29, 0x25, 0x0A, 0x1D, 0x0A, 0x2A, 0x07, 0x4E,
	0x37, 0x2A, 0x05, 0x18, 0x18, 0x07, 0x3C, 0x0F, 0x24, 0x56, 0x07, 0x2E,
	0x7A, 0x3D, 0x2F, 0x45, 0x3D, 0x08, 0x2A, 0x30, 0x1A, 0x3E, 0x03, 0x1D,
	0x02, 0x37, 0x3B, 0x21, 0x5D, 0x17, 0x57, 0x3F, 0x07, 0x2F, 0x58, 0x03,
	0x1F, 0x0E, 0x39, 0x00, 0x09, 0x02, 0x24, 0x1A, 0x38, 0x3A, 0x25, 0x0A,
	0x18, 0x02, 0x28, 0x23, 0x31, 0x1A, 0x10, 0x3D, 0x19, 0x06, 0x0D, 0x59,
	0x1E, 0x27, 0x03, 0x22, 0x24, 0x14, 0x5A, 0x2C, 0x00, 0x0D, 0x3E, 0x23,
	0x0B, 0x2E, 0x11, 0x38, 0x38, 0x73, 0x3C, 0x07, 0x41, 0x00, 0x16, 0x05,
	0x53, 0x05, 0x5E, 0x10, 0x20, 0x0D, 0x5F, 0x28, 0x0A, 0x0A, 0x2A, 0x37,
	0x2A, 0x29, 0x5C, 0x2F, 0x5E, 0x2C, 0x33, 0x1C, 0x07, 0x37, 0x2E, 0x12,
	0x20, 0x35, 0x07, 0x06, 0x07, 0x0B, 0x07, 0x08, 0x22, 0x1A, 0x5A, 0x37,
	0x2D, 0x0C, 0x16, 0x2A, 0x16, 0x0C, 0x19, 0x2B, 0x27, 0x2A, 0x2A, 0x38,
	0x0F, 0x09, 0x08, 0x09, 0x19, 0x00, 0x3E, 0x38, 0x28, 0x07, 0x10, 0x2F,
	0x09, 0x0A, 0x04, 0x25, 0x22, 0x20, 0x0F, 0x2E, 0x23, 0x06, 0x26, 0x05,
	0x07, 0x2A, 0x35, 0x00, 0x25, 0x1C, 0x29, 0x24, 0x06, 0x3E, 0x40, 0x76,
	0x1D, 0x20, 0x0A, 0x3F, 0x07, 0x07, 0x18, 0x36, 0x39, 0x00, 0x00, 0x25,
	0x39, 0x5D, 0x06, 0x1B, 0x18, 0x2A, 0x04, 0x2D, 0x0A, 0x19, 0x25, 0x25,
	0x1A, 0x2F, 0x23, 0x1D, 0x2F, 0x13, 0x2E, 0x38, 0x24, 0x0A, 0x30, 0x28,
	0x4E, 0x36, 0x2E, 0x0F, 0x25, 0x2A, 0x05, 0x32, 0x20, 0x3B, 0x10, 0x1A,
	0x04, 0x04, 0x5E, 0x23, 0x38, 0x53, 0x3A, 0x58, 0x22, 0x45, 0x29, 0x20,
	0x0B, 0x0A, 0x1E, 0x0C, 0x28, 0x2F, 0x29, 0x56, 0x0C, 0x08, 0x58, 0x16,
	0x2A, 0x33, 0x28, 0x24, 0x23, 0x0C, 0x5C, 0x28, 0x16, 0x0C, 0x09, 0x3F,
	0x1A, 0x36, 0x2E, 0x0C, 0x5D, 0x18, 0x0A, 0x39, 0x2C, 0x0A, 0x06, 0x24,
	0x2D, 0x2D, 0x05, 0x17, 0x14, 0x34, 0x3D, 0x1A, 0x74, 0x23, 0x13, 0x3F,
	0x3D, 0x2B, 0x03, 0x22, 0x26, 0x39, 0x1A, 0x18, 0x09, 0x2A, 0x52, 0x03,
	0x06, 0x18, 0x22, 0x3E, 0x00, 0x1A, 0x59, 0x16, 0x04, 0x11, 0x1D, 0x23,
	0x3A, 0x1E, 0x7B, 0x43, 0x55, 0x5D, 0x1B, 0x0D, 0x04, 0x59, 0x3D, 0x3D,
	0x32, 0x25, 0x31, 0x56, 0x2D, 0x74, 0x3A, 0x38, 0x1F, 0x32, 0x18, 0x5B,
	0x31, 0x03, 0x07, 0x15, 0x25, 0x0E, 0x16, 0x06, 0x14, 0x0D, 0x0B, 0x1C,
	0x3F, 0x75, 0x22, 0x08, 0x19, 0x28, 0x0E, 0x2F, 0x30, 0x2F, 0x5E, 0x2A,
	0x07, 0x25, 0x2F, 0x1A, 0x37, 0x08, 0x0D, 0x07, 0x04, 0x0A, 0x2D, 0x03,
	0x02, 0x03, 0x04, 0x06, 0x20, 0x04, 0x3E, 0x0B, 0x21, 0x2B, 0x3C, 0x2E,
	0x15, 0x35, 0x0C, 0x5B, 0x07, 0x04, 0x00, 0x14, 0x5B, 0x2A, 0x2C, 0x54,
	0x35, 0x22, 0x13, 0x27, 0x5D, 0x06, 0x14, 0x02, 0x36, 0x3A, 0x04, 0x09,
	0x27, 0x73, 0x59, 0x15, 0x1C, 0x08, 0x07, 0x0B, 0x38, 0x2D, 0x32, 0x12,
	0x09, 0x28, 0x21, 0x2A, 0x2D, 0x16, 0x1B, 0x09, 0x28, 0x03, 0x25, 0x23,
	0x56, 0x18, 0x00, 0x2D, 0x24, 0x29, 0x2F, 0x0E, 0x2D, 0x51, 0x2C, 0x5F,
	0x17, 0x1B, 0x17, 0x05, 0x2A, 0x11, 0x5D, 0x55, 0x3F, 0x3A, 0x31, 0x36,
	0x10, 0x27, 0x39, 0x2D, 0x1A, 0x31, 0x0B, 0x05, 0x74, 0x39, 0x28, 0x22,
	0x22, 0x21, 0x2E, 0x29, 0x5E, 0x53, 0x72, 0x16, 0x2B, 0x04, 0x58, 0x18,
	0x19, 0x15, 0x2A, 0x2F, 0x2E, 0x25, 0x19, 0x3C, 0x3A, 0x76, 0x1A, 0x06,
	0x3B, 0x05, 0x0F, 0x38, 0x38, 0x1F, 0x00, 0x1A, 0x39, 0x23, 0x45, 0x53,
	0x2D, 0x23, 0x05, 0x18, 0x09, 0x34, 0x09, 0x04, 0x1E, 0x07, 0x26, 0x0B,
	0x03, 0x18, 0x00, 0x27, 0x02, 0x14, 0x21, 0x2D, 0x14, 0x1B, 0x2C, 0x29,
	0x1C, 0x1A, 0x1C, 0x30, 0x16, 0x5D, 0x0D, 0x0F, 0x00, 0x58, 0x38, 0x27,
	0x3C, 0x30, 0x2C, 0x31, 0x1B, 0x26, 0x50, 0x01, 0x07, 0x33, 0x28, 0x0C,
	0x02, 0x19, 0x06, 0x01, 0x0D, 0x1F, 0x2F, 0x2F, 0x5C, 0x59, 0x5B, 0x28,
	0x29, 0x03, 0x16, 0x04, 0x40, 0x1B, 0x39, 0x0A, 0x3E, 0x3E, 0x07, 0x1A,
	0x24, 0x22, 0x5C, 0x75, 0x1C, 0x27, 0x24, 0x29, 0x35, 0x3F, 0x09, 0x07,
	0x07, 0x13, 0x5E, 0x15, 0x59, 0x22, 0x33, 0x28, 0x20, 0x0D, 0x59, 0x2B,
	0x20, 0x24, 0x29, 0x09, 0x70, 0x20, 0x29, 0x2B, 0x1C, 0x11, 0x2F, 0x32,
	0x37, 0x3A, 0x2F, 0x14, 0x2B, 0x16, 0x28, 0x16, 0x2B, 0x2A, 0x3E, 0x21,
	0x29, 0x39, 0x58, 0x38, 0x09, 0x72, 0x14, 0x4A, 0x00, 0x33, 0x0B, 0x59,
	0x50, 0x36, 0x3A, 0x04, 0x54, 0x32, 0x00, 0x02, 0x24, 0x2F, 0x4E, 0x37,
	0x3D, 0x7A, 0x0D, 0x35, 0x3D, 0x39, 0x0D, 0x21, 0x54, 0x36, 0x3C, 0x25,
	0x03, 0x52, 0x36, 0x44, 0x05, 0x01, 0x0C, 0x2F, 0x2E, 0x1B, 0x05, 0x53,
	0x2F, 0x04, 0x2C, 0x07, 0x4E, 0x24, 0x18, 0x03, 0x5E, 0x54, 0x41, 0x18,
	0x17, 0x3F, 0x52, 0x01, 0x38, 0x77, 0x22, 0x24, 0x0B, 0x52, 0x32, 0x28,
	0x22, 0x09, 0x09, 0x74, 0x28, 0x1B, 0x21, 0x1B, 0x0A, 0x00, 0x0F, 0x0D,
	0x0A, 0x73, 0x35, 0x08, 0x2A, 0x1E, 0x77, 0x38, 0x0C, 0x26, 0x0C, 0x26,
	0x01, 0x2C, 0x03, 0x2A, 0x37, 0x3F, 0x58, 0x2A, 0x07, 0x3A, 0x54, 0x2F,
	0x5E, 0x18, 0x1A, 0x47, 0x2A, 0x3C, 0x58, 0x16, 0x01, 0x22, 0x39, 0x03,
	0x37, 0x1A, 0x55, 0x03, 0x29, 0x13, 0x1F, 0x4E, 0x2A, 0x38, 0x70, 0x29,
	0x32, 0x59, 0x11, 0x14, 0x03, 0x2D, 0x39, 0x26, 0x0D, 0x1C, 0x06, 0x04,
	0x09, 0x20, 0x03, 0x17, 0x18, 0x2C, 0x35, 0x3B, 0x05, 0x03, 0x06, 0x33,
	0x2B, 0x0F, 0x04, 0x25, 0x2C, 0x0A, 0x26, 0x2A, 0x25, 0x2D, 0x0F, 0x0F,
	0x05, 0x52, 0x34, 0x21, 0x13, 0x34, 0x32, 0x0D, 0x3E, 0x23, 0x37, 0x2A,
	0x03, 0x08, 0x4A, 0x36, 0x2D, 0x0E, 0x5B, 0x27, 0x37, 0x28, 0x69, 0x2F,
	0x51, 0x3A, 0x3C, 0x25, 0x5B, 0x13, 0x59, 0x27, 0x2B, 0x0E, 0x0E, 0x08,
	0x39, 0x10, 0x22, 0x16, 0x59, 0x3F, 0x0F, 0x3C, 0x07, 0x01, 0x25, 0x14,
	0x19, 0x32, 0x29, 0x24, 0x69, 0x03, 0x52, 0x37, 0x2D, 0x38, 0x3F, 0x4A,
	0x57, 0x18, 0x30, 0x0A, 0x2B, 0x0D, 0x3B, 0x30, 0x2F, 0x2D, 0x23, 0x33,
	0x17, 0x00, 0x19, 0x36, 0x3F, 0x30, 0x5E, 0x52, 0x2B, 0x06, 0x7A, 0x18,
	0x29, 0x14, 0x2A, 0x71, 0x2E, 0x07, 0x5D, 0x5C, 0x0C, 0x5E, 0x4A, 0x2C,
	0x28, 0x2D, 0x5C, 0x12, 0x20, 0x1C, 0x11, 0x5A, 0x39, 0x16, 0x01, 0x25,
	0x26, 0x53, 0x5D, 0x1D, 0x71, 0x47, 0x04, 0x20, 0x28, 0x04, 0x0B, 0x04,
	0x0A, 0x31, 0x32, 0x3D, 0x54, 0x38, 0x2F, 0x70, 0x5D, 0x31, 0x18, 0x44,
	0x17, 0x2B, 0x23, 0x36, 0x21, 0x33, 0x58, 0x0E, 0x5E, 0x0A, 0x20, 0x54,
	0x57, 0x39, 0x3C, 0x1B, 0x3C, 0x34, 0x3C, 0x23, 0x0E, 0x39, 0x09, 0x0D,
	0x01, 0x3B, 0x1E, 0x31, 0x39, 0x3E, 0x18, 0x39, 0x4E, 0x09, 0x39, 0x21,
	0x5A, 0x53, 0x2B, 0x53, 0x0E, 0x3B, 0x0F, 0x14, 0x1B, 0x32, 0x34, 0x22,
	0x1C, 0x1C, 0x0E, 0x25, 0x13, 0x5E, 0x1C, 0x21, 0x1A, 0x16, 0x0A, 0x40,
	0x38, 0x5E, 0x28, 0x05, 0x5C, 0x23, 0x43, 0x28, 0x00, 0x5D, 0x28, 0x3E,
	0x32, 0x03, 0x1D, 0x29, 0x0A, 0x08, 0x39, 0x39, 0x27, 0x05, 0x53, 0x04,
	0x2F, 0x15, 0x58, 0x30, 0x0F, 0x07, 0x17, 0x2A, 0x29, 0x03, 0x40, 0x01,
	0x2F, 0x30, 0x1C, 0x1E, 0x6D, 0x59, 0x26, 0x23, 0x1B, 0x74, 0x2A, 0x18,
	0x2C, 0x31, 0x08, 0x2A, 0x4E, 0x3A, 0x07, 0x18, 0x29, 0x56, 0x16, 0x13,
	0x01, 0x3F, 0x32, 0x14, 0x40, 0x14, 0x5C, 0x18, 0x18, 0x2A, 0x75, 0x5E,
	0x28, 0x5E, 0x07, 0x17, 0x29, 0x59, 0x16, 0x3F, 0x07, 0x18, 0x16, 0x39,
	0x2F, 0x06, 0x0B, 0x03, 0x2D, 0x39, 0x32, 0x2D, 0x0D, 0x16, 0x24, 0x34,
	0x25, 0x27, 0x5E, 0x2A, 0x15, 0x34, 0x10, 0x2C, 0x3A, 0x04, 0x58, 0x13,
	0x2A, 0x20, 0x03, 0x5A, 0x03, 0x5F, 0x5A, 0x09, 0x5D, 0x31, 0x05, 0x28,
	0x0F, 0x0B, 0x23, 0x41, 0x52, 0x3A, 0x5A, 0x27, 0x23, 0x2A, 0x06, 0x0A,
	0x20, 0x2A, 0x12, 0x36, 0x23, 0x2B, 0x3A, 0x3B, 0x01, 0x3E, 0x52, 0x04,
	0x03, 0x77, 0x15, 0x50, 0x0A, 0x13, 0x09, 0x5D, 0x53, 0x00, 0x3F, 0x34,
	0x18, 0x52, 0x09, 0x0C, 0x0C, 0x0D, 0x2A, 0x5E, 0x06, 0x07, 0x04, 0x39,
	0x57, 0x3B, 0x36, 0x5C, 0x4E, 0x06, 0x21, 0x1B, 0x03, 0x07, 0x29, 0x44,
	0x16, 0x1B, 0x23, 0x5A, 0x33, 0x3A, 0x09, 0x16, 0x17, 0x19, 0x06, 0x0A,
	0x11, 0x2D, 0x29, 0x76, 0x24, 0x16, 0x04, 0x1F, 0x33, 0x20, 0x38, 0x09,
	0x53, 0x16, 0x39, 0x26, 0x3E, 0x22, 0x73, 0x47, 0x0A, 0x0F, 0x01, 0x34,
	0x5F, 0x57, 0x07, 0x20, 0x2D, 0x2D, 0x11, 0x2B, 0x27, 0x73, 0x2F, 0x57,
	0x3C, 0x44, 0x1B, 0x2F, 0x07, 0x14, 0x01, 0x31, 0x08, 0x23, 0x1B, 0x0D,
	0x29, 0x2A, 0x18, 0x36, 0x01, 0x38, 0x1F, 0x0D, 0x06, 0x33, 0x11, 0x07,
	0x57, 0x3C, 0x2E, 0x26, 0x1C, 0x35, 0x57, 0x38, 0x10, 0x25, 0x24, 0x27,
	0x5D, 0x11, 0x1D, 0x55, 0x00, 0x1C, 0x03, 0x26, 0x33, 0x34, 0x29, 0x0A,
	0x21, 0x03, 0x17, 0x0E, 0x0E, 0x09, 0x57, 0x3D, 0x01, 0x1B, 0x3E, 0x09,
	0x14, 0x29, 0x35, 0x2F, 0x59, 0x5C, 0x2A, 0x72, 0x29, 0x52, 0x00, 0x29,
	0x0F, 0x0D, 0x08, 0x19, 0x3C, 0x18, 0x3A, 0x36, 0x2F, 0x3F, 0x26, 0x29,
	0x30, 0x1F, 0x52, 0x2F, 0x29, 0x32, 0x17, 0x07, 0x06, 0x08, 0x0F, 0x09,
	0x5D, 0x1B, 0x5D, 0x59, 0x5D, 0x18, 0x30, 0x2D, 0x10, 0x5E, 0x1F, 0x76,
	0x5D, 0x38, 0x2D, 0x33, 0x01, 0x07, 0x02, 0x05, 0x27, 0x17, 0x39, 0x08,
	0x3A, 0x3E, 0x17, 0x05, 0x38, 0x3D, 0x1C, 0x77, 0x07, 0x24, 0x03, 0x29,
	0x04, 0x26, 0x02, 0x19, 0x1B, 0x12, 0x28, 0x32, 0x5C, 0x29, 0x2D, 0x03,
	0x0C, 0x3D, 0x29, 0x18, 0x05, 0x23, 0x25, 0x09, 0x0B, 0x3B, 0x39, 0x2C,
	0x2E, 0x35, 0x15, 0x17, 0x28, 0x11, 0x0F, 0x23, 0x16, 0x2F, 0x03, 0x03,
	0x1C, 0x20, 0x3E, 0x00, 0x77, 0x0F, 0x2A, 0x09, 0x29, 0x2A, 0x05, 0x18,
	0x01, 0x53, 0x09, 0x3D, 0x10, 0x1D, 0x2D, 0x17, 0x16, 0x26, 0x2B, 0x26,
	0x1B, 0x43, 0x57, 0x06, 0x07, 0x31, 0x3C, 0x28, 0x26, 0x28, 0x17, 0x1D,
	0x17, 0x0F, 0x3A, 0x0C, 0x04, 0x19, 0x0A, 0x2F, 0x0B, 0x16, 0x4E, 0x2C,
	0x21, 0x76, 0x19, 0x2B, 0x57, 0x52, 0x18, 0x55, 0x30, 0x5F, 0x22, 0x07,
	0x3A, 0x2E, 0x0F, 0x5B, 0x04, 0x1C, 0x30, 0x09, 0x27, 0x18, 0x23, 0x28,
	0x02, 0x52, 0x75, 0x47, 0x20, 0x01, 0x0E, 0x71, 0x3D, 0x2F, 0x26, 0x04,
	0x04, 0x22, 0x36, 0x2B, 0x0E, 0x00, 0x04, 0x00, 0x2A, 0x5B, 0x00, 0x09,
	0x53, 0x3E, 0x25, 0x2D, 0x04, 0x51, 0x58, 0x01, 0x1A, 0x0B, 0x00, 0x41,
	0x38, 0x17, 0x24, 0x31, 0x14, 0x20, 0x12, 0x25, 0x30, 0x16, 0x0D, 0x2F,
	0x0B, 0x0F, 0x45, 0x2E, 0x06, 0x38, 0x52, 0x3F, 0x1D, 0x76, 0x3D, 0x00,
	0x24, 0x3C, 0x70, 0x5A, 0x30, 0x1C, 0x0E, 0x15, 0x3A, 0x38, 0x07, 0x0D,
	0x05, 0x21, 0x53, 0x5E, 0x3A, 0x3A, 0x04, 0x55, 0x2B, 0x3C, 0x10, 0x38,
	0x23, 0x3B, 0x21, 0x14, 0x2A, 0x0E, 0x04, 0x25, 0x0B, 0x20, 0x59, 0x3C,
	0x26, 0x3A, 0x0F, 0x30, 0x1F, 0x5F, 0x73, 0x1D, 0x23, 0x5B, 0x5D, 0x71,
	0x00, 0x2C, 0x1A, 0x0D, 0x0D, 0x35, 0x1B, 0x3C, 0x2F, 0x2C, 0x09, 0x59,
	0x09, 0x1A, 0x38, 0x54, 0x20, 0x3A, 0x04, 0x09, 0x15, 0x04, 0x3F, 0x32,
	0x29, 0x0E, 0x16, 0x5F, 0x2C, 0x14, 0x29, 0x2E, 0x2B, 0x58, 0x26, 0x27,
	0x08, 0x39, 0x23, 0x04, 0x21, 0x26, 0x3B, 0x1C, 0x11, 0x0B, 0x0F, 0x3C,
	0x1C, 0x7B, 0x2E, 0x52, 0x2F, 0x0D, 0x14, 0x5A, 0x58, 0x27, 0x22, 0x0E,
	0x03, 0x08, 0x17, 0x1A, 0x17, 0x5D, 0x39, 0x1C, 0x32, 0x05, 0x35, 0x15,
	0x01, 0x5F, 0x30, 0x3D, 0x30, 0x45, 0x3C, 0x73, 0x3D, 0x56, 0x3A, 0x09,
	0x37, 0x25, 0x08, 0x09, 0x23, 0x27, 0x0F, 0x13, 0x5A, 0x27, 0x73, 0x3B,
	0x54, 0x3B, 0x19, 0x0B, 0x23, 0x3B, 0x22, 0x0C, 0x33, 0x1D, 0x55, 0x3B,
	0x1A, 0x2D, 0x29, 0x2D, 0x26, 0x3D, 0x20, 0x5D, 0x33, 0x23, 0x2D, 0x10,
	0x3A, 0x38, 0x06, 0x3C, 0x0D, 0x2E, 0x0D, 0x2B, 0x1E, 0x14, 0x02, 0x20,
	0x3A, 0x1C, 0x26, 0x05, 0x19, 0x01, 0x59, 0x11, 0x1B, 0x09, 0x1D, 0x01,
	0x21, 0x1E, 0x2C, 0x02, 0x01, 0x00, 0x18, 0x0E, 0x18, 0x2A, 0x0E, 0x21,
	0x07, 0x18, 0x5B, 0x3A, 0x23, 0x0D, 0x0D, 0x1E, 0x3A, 0x39, 0x29, 0x07,
	0x24, 0x2A, 0x2D, 0x31, 0x08, 0x09, 0x17, 0x5D, 0x57, 0x2B, 0x02, 0x30,
	0x43, 0x2A, 0x2B, 0x32, 0x3B, 0x2E, 0x08, 0x27, 0x1D, 0x38, 0x19, 0x0B,
	0x1C, 0x00, 0x01, 0x28, 0x58, 0x24, 0x5B, 0x37, 0x2B, 0x06, 0x27, 0x27,
	0x1B, 0x1D, 0x27, 0x29, 0x28, 0x15, 0x58, 0x26, 0x22, 0x53, 0x0E, 0x1E,
	0x11, 0x0B, 0x01, 0x00, 0x54, 0x2A, 0x2C, 0x5A, 0x0A, 0x0F, 0x2A, 0x59,
	0x27, 0x76, 0x02, 0x52, 0x3A, 0x19, 0x10, 0x1E, 0x12, 0x38, 0x24, 0x06,
	0x2F, 0x3B, 0x3E, 0x2A, 0x34, 0x5D, 0x16, 0x3C, 0x09, 0x01, 0x0B, 0x07,
	0x56, 0x28, 0x7A, 0x5F, 0x20, 0x14, 0x0A, 0x11, 0x27, 0x0C, 0x17, 0x00,
	0x1A, 0x1D, 0x52, 0x16, 0x21, 0x09, 0x55, 0x37, 0x2B, 0x39, 0x34, 0x3A,
	0x55, 0x08, 0x18, 0x0E, 0x3D, 0x32, 0x0A, 0x1A, 0x06, 0x09, 0x18, 0x27,
	0x3D, 0x3B, 0x20, 0x0B, 0x2D, 0x59, 0x01, 0x54, 0x03, 0x3B, 0x0E, 0x7A,
	0x02, 0x25, 0x0B, 0x3F, 0x1B, 0x34, 0x1B, 0x3E, 0x01, 0x2C, 0x0B, 0x50,
	0x23, 0x1B, 0x75, 0x5D, 0x20, 0x58, 0x06, 0x0F, 0x06, 0x2D, 0x0A, 0x0A,
	0x23, 0x23, 0x16, 0x2C, 0x3F, 0x07, 0x19, 0x03, 0x2A, 0x06, 0x69, 0x21,
	0x30, 0x3A, 0x58, 0x3A, 0x3A, 0x39, 0x29, 0x23, 0x2D, 0x26, 0x2B, 0x3F,
	0x0E, 0x38, 0x3E, 0x33, 0x5E, 0x2E, 0x35, 0x2B, 0x00, 0x09, 0x13, 0x25,
	0x28, 0x26, 0x19, 0x02, 0x3A, 0x36, 0x13, 0x1D, 0x2D, 0x25, 0x3B, 0x35,
	0x5B, 0x1A, 0x36, 0x2E, 0x2E, 0x18, 0x5C, 0x76, 0x1C, 0x02, 0x3F, 0x1B,
	0x0D, 0x39, 0x51, 0x04, 0x5C, 0x2E, 0x1C, 0x10, 0x38, 0x1B, 0x1B, 0x5E,
	0x00, 0x1D, 0x28, 0x18, 0x5B, 0x50, 0x05, 0x06, 0x0F, 0x1D, 0x29, 0x0F,
	0x5D, 0x13, 0x2A, 0x30, 0x1A, 0x19, 0x27, 0x28, 0x07, 0x29, 0x1A, 0x32,
	0x3B, 0x53, 0x57, 0x39, 0x72, 0x23, 0x06, 0x29, 0x29, 0x0C, 0x38, 0x06,
	0x24, 0x3E, 0x28, 0x5B, 0x07, 0x1C, 0x20, 0x1B, 0x3B, 0x2D, 0x07, 0x38,
	0x17, 0x2A, 0x17, 0x27, 0x44, 0x34, 0x20, 0x16, 0x1B, 0x5B, 0x35, 0x01,
	0x31, 0x08, 0x0A, 0x0C, 0x3D, 0x27, 0x22, 0x53, 0x2B, 0x00, 0x23, 0x3C,
	0x38, 0x06, 0x16, 0x25, 0x3D, 0x22, 0x07, 0x2E, 0x50, 0x25, 0x2A, 0x2D,
	0x23, 0x17, 0x09, 0x58, 0x0A, 0x04, 0x13, 0x1E, 0x38, 0x25, 0x2F, 0x3B,
	0x3F, 0x04, 0x20, 0x16, 0x20, 0x02, 0x21, 0x06, 0x16, 0x2A, 0x06, 0x23,
	0x25, 0x0B, 0x33, 0x5E, 0x2C, 0x09, 0x2E, 0x37, 0x23, 0x3C, 0x03, 0x0D,
	0x33, 0x04, 0x3B, 0x72, 0x3D, 0x02, 0x5C, 0x21, 0x0B, 0x35, 0x34, 0x45,
	0x1A, 0x07, 0x00, 0x23, 0x41, 0x0F, 0x1A, 0x25, 0x24, 0x1C, 0x5E, 0x1A,
	0x28, 0x0D, 0x5A, 0x3A, 0x14, 0x54, 0x12, 0x0F, 0x28, 0x0C, 0x07, 0x34,
	0x5F, 0x00, 0x71, 0x29, 0x28, 0x3A, 0x07, 0x07, 0x00, 0x35, 0x36, 0x28,
	0x74, 0x38, 0x02, 0x06, 0x58, 0x32, 0x58, 0x20, 0x3E, 0x0A, 0x01, 0x15,
	0x0C, 0x41, 0x27, 0x18, 0x0B, 0x3B, 0x57, 0x0F, 0x08, 0x5F, 0x51, 0x29,
	0x2F, 0x05, 0x35, 0x0A, 0x34, 0x5F, 0x0C, 0x54, 0x06, 0x28, 0x04, 0x0D,
	0x1A, 0x55, 0x0C, 0x39, 0x12, 0x0A, 0x52, 0x56, 0x2A, 0x37, 0x00, 0x28,
	0x0B, 0x20, 0x04, 0x25, 0x03, 0x45, 0x3C, 0x11, 0x36, 0x09, 0x19, 0x22,
	0x09, 0x03, 0x51, 0x1F, 0x1F, 0x12, 0x0F, 0x2D, 0x00, 0x19, 0x73, 0x38,
	0x11, 0x3E, 0x08, 0x07, 0x55, 0x25, 0x06, 0x25, 0x2F, 0x1B, 0x0A, 0x5D,
	0x2D, 0x2C, 0x02, 0x2E, 0x2F, 0x3D, 0x74, 0x2E, 0x0F, 0x5C, 0x0F, 0x24,
	0x2B, 0x27, 0x20, 0x5D, 0x01, 0x19, 0x33, 0x25, 0x0E, 0x05, 0x0A, 0x22,
	0x1E, 0x38, 0x14, 0x3C, 0x2F, 0x3C, 0x3A, 0x20, 0x1C, 0x4E, 0x2A, 0x24,
	0x0A, 0x2D, 0x14, 0x57, 0x53, 0x12, 0x1B, 0x0D, 0x1C, 0x3F, 0x13, 0x2D,
	0x04, 0x1F, 0x00, 0x25, 0x3A, 0x14, 0x04, 0x08, 0x76, 0x0B, 0x07, 0x56,
	0x3D, 0x09, 0x2A, 0x2C, 0x20, 0x1A, 0x09, 0x07, 0x35, 0x37, 0x26, 0x70,
	0x29, 0x58, 0x59, 0x01, 0x71, 0x39, 0x34, 0x36, 0x3B, 0x28, 0x27, 0x4E,
	0x3F, 0x13, 0x24, 0x09, 0x2E, 0x34, 0x44, 0x17, 0x04, 0x37, 0x26, 0x58,
	0x12, 0x3D, 0x2D, 0x3E, 0x19, 0x72, 0x18, 0x29, 0x58, 0x58, 0x14, 0x03,
	0x30, 0x22, 0x02, 0x2D, 0x22, 0x4A, 0x1E, 0x27, 0x3A, 0x2E, 0x2F, 0x36,
	0x3B, 0x14, 0x06, 0x03, 0x26, 0x5D, 0x25, 0x27, 0x0B, 0x5B, 0x29, 0x37,
	0x28, 0x0F, 0x3F, 0x00, 0x15, 0x01, 0x0A, 0x04, 0x59, 0x23, 0x55, 0x33,
	0x27, 0x07, 0x2F, 0x55, 0x31, 0x2F, 0x3D, 0x07, 0x02, 0x59, 0x09, 0x3C,
	0x21, 0x1D, 0x4E, 0x5E, 0x06, 0x69, 0x58, 0x17, 0x1D, 0x00, 0x14, 0x3C,
	0x0C, 0x00, 0x3E, 0x75, 0x1F, 0x08, 0x5D, 0x1D, 0x3B, 0x24, 0x00, 0x58,
	0x3B, 0x04, 0x1A, 0x0D, 0x14, 0x1F, 0x2F, 0x5E, 0x02, 0x09, 0x2C, 0x7B,
	0x0F, 0x34, 0x36, 0x3C, 0x74, 0x2F, 0x2D, 0x3F, 0x25, 0x14, 0x5E, 0x18,
	0x26, 0x00, 0x00, 0x07, 0x0B, 0x34, 0x5D, 0x17, 0x5A, 0x02, 0x24, 0x21,
	0x17, 0x3E, 0x14, 0x37, 0x53, 0x07, 0x1E, 0x07, 0x08, 0x5E, 0x16, 0x26,
	0x54, 0x26, 0x07, 0x1B, 0x03, 0x18, 0x25, 0x2E, 0x03, 0x5D, 0x29, 0x5C,
	0x0A, 0x2E, 0x5E, 0x18, 0x5F, 0x5E, 0x26, 0x5B, 0x2F, 0x2D, 0x1B, 0x20,
	0x3A, 0x34, 0x03, 0x39, 0x00, 0x2F, 0x00, 0x2B, 0x06, 0x0F, 0x0B, 0x2C,
	0x5D, 0x07, 0x26, 0x5E, 0x06, 0x45, 0x29, 0x03, 0x2D, 0x59, 0x2C, 0x3D,
	0x75, 0x5E, 0x59, 0x01, 0x06, 0x07, 0x34, 0x36, 0x3F, 0x23, 0x1B, 0x0D,
	0x2F, 0x26, 0x31, 0x15, 0x43, 0x0E, 0x1E, 0x0D, 0x11, 0x24, 0x57, 0x39,
	0x3E, 0x01, 0x07, 0x52, 0x5E, 0x33, 0x3B, 0x3C, 0x0F, 0x2D, 0x31, 0x0C,
	0x23, 0x30, 0x1C, 0x1F, 0x74, 0x14, 0x25, 0x59, 0x3F, 0x12, 0x3D, 0x28,
	0x14, 0x39, 0x0F, 0x23, 0x09, 0x03, 0x5A, 0x35, 0x24, 0x0E, 0x39, 0x1C,
	0x05, 0x25, 0x15, 0x29, 0x06, 0x2B, 0x04, 0x05, 0x23, 0x39, 0x30, 0x54,
	0x51, 0x28, 0x0C, 0x30, 0x28, 0x0E, 0x20, 0x3F, 0x31, 0x3D, 0x36, 0x19,
	0x0E, 0x06, 0x3F, 0x04, 0x3B, 0x13, 0x7A, 0x06, 0x17, 0x3B, 0x5E, 0x2B,
	0x18, 0x28, 0x08, 0x2A, 0x33, 0x2D, 0x51, 0x0F, 0x5F, 0x01, 0x29, 0x06,
	0x0A, 0x39, 0x15, 0x21, 0x2A, 0x1F, 0x0E, 0x2F, 0x27, 0x23, 0x22, 0x19,
	0x12, 0x03, 0x26, 0x24, 0x28, 0x14, 0x24, 0x02, 0x0B, 0x0A, 0x11, 0x24,
	0x22, 0x2B, 0x1B, 0x13, 0x23, 0x12, 0x3D, 0x07, 0x11, 0x26, 0x0D, 0x34,
	0x38, 0x24, 0x2F, 0x2D, 0x02, 0x0E, 0x0E, 0x00, 0x27, 0x37, 0x52, 0x13,
	0x3F, 0x30, 0x1F, 0x2C, 0x32, 0x5F, 0x10, 0x06, 0x39, 0x76, 0x15, 0x52,
	0x1C, 0x3D, 0x05, 0x29, 0x19, 0x2F, 0x32, 0x09, 0x18, 0x12, 0x07, 0x2D,
	0x35, 0x2A, 0x4A, 0x3E, 0x06, 0x06, 0x14, 0x57, 0x19, 0x58, 0x75, 0x3A,
	0x24, 0x17, 0x38, 0x06, 0x22, 0x56, 0x5D, 0x2A, 0x01, 0x28, 0x0D, 0x1F,
	0x32, 0x17, 0x3D, 0x38, 0x57, 0x27, 0x10, 0x35, 0x29, 0x39, 0x22, 0x09,
	0x2F, 0x24, 0x21, 0x1C, 0x2B, 0x1A, 0x2D, 0x36, 0x5E, 0x06, 0x1E, 0x55,
	0x36, 0x58, 0x01, 0x0F, 0x14, 0x2D, 0x5C, 0x0A, 0x25, 0x07, 0x3A, 0x13,
	0x20, 0x15, 0x0E, 0x09, 0x04, 0x15, 0x5A, 0x54, 0x04, 0x02, 0x13, 0x0E,
	0x16, 0x3A, 0x01, 0x2E, 0x5D, 0x24, 0x03, 0x20, 0x26, 0x59, 0x55, 0x5E,
	0x2E, 0x3A, 0x3F, 0x08, 0x38, 0x1A, 0x03, 0x03, 0x2C, 0x28, 0x18, 0x0E,
	0x25, 0x27, 0x3F, 0x23, 0x7B, 0x24, 0x30, 0x04, 0x3A, 0x16, 0x54, 0x51,
	0x57, 0x5D, 0x1A, 0x01, 0x31, 0x3D, 0x20, 0x14, 0x3D, 0x36, 0x21, 0x28,
	0x10, 0x0A, 0x30, 0x27, 0x18, 0x2D, 0x09, 0x11, 0x05, 0x0F, 0x28, 0x27,
	0x26, 0x01, 0x0C, 0x0B, 0x0E, 0x58, 0x5C, 0x24, 0x32, 0x18, 0x0E, 0x3E,
	0x28, 0x2E, 0x22, 0x36, 0x28, 0x27, 0x20, 0x1E, 0x24, 0x0F, 0x07, 0x27,
	0x08, 0x34, 0x39, 0x1D, 0x70, 0x1B, 0x32, 0x37, 0x3D, 0x2C, 0x1D, 0x3B,
	0x03, 0x20, 0x7B, 0x38, 0x00, 0x2A, 0x26, 0x34, 0x07, 0x0B, 0x20, 0x58,
	0x15, 0x19, 0x0D, 0x0B, 0x1E, 0x15, 0x43, 0x0C, 0x27, 0x08, 0x09, 0x24,
	0x22, 0x3C, 0x58, 0x2A, 0x0E, 0x2B, 0x5B, 0x3C, 0x36, 0x0B, 0x0D, 0x24,
	0x5D, 0x6D, 0x21, 0x2F, 0x1F, 0x23, 0x72, 0x21, 0x38, 0x3E, 0x18, 0x71,
	0x15, 0x20, 0x1B, 0x5B, 0x10, 0x0B, 0x39, 0x39, 0x3E, 0x28, 0x0F, 0x53,
	0x2B, 0x24, 0x31, 0x24, 0x13, 0x37, 0x3D, 0x11, 0x27, 0x37, 0x16, 0x26,
	0x2D, 0x3F, 0x55, 0x28, 0x2E, 0x17, 0x2E, 0x03, 0x2B, 0x3C, 0x15, 0x2F,
	0x33, 0x2F, 0x18, 0x20, 0x15, 0x2B, 0x1C, 0x3F, 0x0D, 0x47, 0x29, 0x41,
	0x07, 0x2F, 0x05, 0x2A, 0x0F, 0x06, 0x2F, 0x06, 0x27, 0x1A, 0x23, 0x14,
	0x23, 0x14, 0x1E, 0x5B, 0x2F, 0x5D, 0x0D, 0x22, 0x01, 0x15, 0x1F, 0x06,
	0x06, 0x23, 0x25, 0x18, 0x05, 0x3D, 0x3F, 0x32, 0x0B, 0x4E, 0x1B, 0x18,
	0x04, 0x23, 0x34, 0x39, 0x3B, 0x29, 0x3D, 0x37, 0x5F, 0x31, 0x07, 0x19,
	0x07, 0x3F, 0x08, 0x1B, 0x3A, 0x34, 0x5E, 0x20, 0x0C, 0x47, 0x2E, 0x2C,
	0x0A, 0x2C, 0x08, 0x00, 0x29, 0x0E, 0x28, 0x0B, 0x4E, 0x5E, 0x5E, 0x11,
	0x2A, 0x0B, 0x38, 0x13, 0x05, 0x55, 0x20, 0x58, 0x3E, 0x28, 0x15, 0x25,
	0x16, 0x1C, 0x30, 0x26, 0x07, 0x06, 0x29, 0x01, 0x27, 0x27, 0x3A, 0x2F,
	0x76, 0x0E, 0x20, 0x2A, 0x08, 0x21, 0x20, 0x13, 0x5B, 0x3C, 0x31, 0x3E,
	0x30, 0x2A, 0x5D, 0x05, 0x21, 0x35, 0x2C, 0x26, 0x2C, 0x18, 0x20, 0x2D,
	0x04, 0x14, 0x00, 0x18, 0x29, 0x00, 0x32, 0x47, 0x2A, 0x38, 0x3F, 0x13,
	0x39, 0x24, 0x0F, 0x0A, 0x11, 0x07, 0x2D, 0x28, 0x1E, 0x29, 0x3C, 0x29,
	0x01, 0x00, 0x04, 0x5F, 0x2B, 0x3C, 0x0A, 0x15, 0x1E, 0x18, 0x06, 0x2F,
	0x2E, 0x15, 0x09, 0x2A, 0x3C, 0x31, 0x1A, 0x55, 0x3D, 0x2E, 0x32, 0x1A,
	0x0A, 0x24, 0x3C, 0x71, 0x25, 0x04, 0x5F, 0x1C, 0x12, 0x3A, 0x2D, 0x59,
	0x1C, 0x07, 0x23, 0x08, 0x05, 0x2F, 0x23, 0x07, 0x18, 0x2F, 0x2F, 0x21,
	0x18, 0x28, 0x2F, 0x3A, 0x26, 0x3D, 0x07, 0x25, 0x04, 0x01, 0x07, 0x2A,
	0x06, 0x06, 0x2F, 0x3E, 0x2A, 0x07, 0x29, 0x13, 0x25, 0x0D, 0x29, 0x53,
	0x13, 0x2D, 0x37, 0x29, 0x1F, 0x08, 0x1D, 0x36, 0x23, 0x2F, 0x75, 0x05,
	0x34, 0x2A, 0x06, 0x73, 0x26, 0x29, 0x20, 0x3E, 0x03, 0x0F, 0x10, 0x38,
	0x24, 0x69, 0x21, 0x0B, 0x41, 0x5D, 0x2B, 0x0F, 0x3B, 0x3A, 0x18, 0x13,
	0x54, 0x4A, 0x5A, 0x0C, 0x11, 0x1E, 0x36, 0x5E, 0x3D, 0x10, 0x21, 0x4A,
	0x0C, 0x3D, 0x12, 0x20, 0x28, 0x3A, 0x18, 0x24, 0x0F, 0x05, 0x5E, 0x0E,
	0x7B, 0x08, 0x37, 0x0D, 0x21, 0x00, 0x3E, 0x30, 0x38, 0x3C, 0x07, 0x15,
	0x4A, 0x2B, 0x59, 0x70, 0x3D, 0x52, 0x14, 0x00, 0x07, 0x2F, 0x0E, 0x1B,
	0x3C, 0x11, 0x39, 0x11, 0x1F, 0x3D, 0x7B, 0x5E, 0x37, 0x25, 0x06, 0x77,
	0x03, 0x51, 0x1C, 0x25, 0x2C, 0x0D, 0x15, 0x05, 0x39, 0x13, 0x03, 0x35,
	0x5D, 0x3A, 0x76, 0x22, 0x30, 0x1F, 0x28, 0x08, 0x20, 0x28, 0x36, 0x44,
	0x2D, 0x04, 0x03, 0x20, 0x05, 0x15, 0x1C, 0x33, 0x25, 0x5D, 0x69, 0x2A,
	0x05, 0x5F, 0x0D, 0x0D, 0x2E, 0x11, 0x04, 0x5D, 0x38, 0x05, 0x39, 0x28,
	0x2D, 0x7A, 0x00, 0x35, 0x3D, 0x07, 0x72, 0x1B, 0x56, 0x37, 0x3B, 0x33,
	0x23, 0x34, 0x3D, 0x40, 0x3A, 0x04, 0x32, 0x02, 0x32, 0x0E, 0x5C, 0x38,
	0x21, 0x21, 0x71, 0x19, 0x53, 0x02, 0x26, 0x29, 0x5D, 0x2C, 0x56, 0x3D,
	0x1A, 0x0A, 0x2C, 0x58, 0x52, 0x0E, 0x22, 0x1B, 0x36, 0x1D, 0x16, 0x0A,
	0x2C, 0x09, 0x1E, 0x08, 0x0D, 0x3B, 0x08, 0x53, 0x11, 0x2F, 0x11, 0x3A,
	0x5A, 0x73, 0x08, 0x51, 0x1E, 0x3C, 0x10, 0x05, 0x0D, 0x14, 0x11, 0x38,
	0x43, 0x0E, 0x0B, 0x3E, 0x0A, 0x29, 0x2D, 0x09, 0x32, 0x25, 0x5A, 0x50,
	0x37, 0x3F, 0x32, 0x04, 0x4A, 0x06, 0x40, 0x37, 0x0B, 0x09, 0x28, 0x00,
	0x0A, 0x21, 0x20, 0x1D, 0x12, 0x26, 0x20, 0x27, 0x08, 0x5B, 0x24, 0x20,
	0x02, 0x59, 0x40, 0x2B, 0x1C, 0x38, 0x3A, 0x5D, 0x30, 0x0E, 0x19, 0x1C,
	0x58, 0x1B, 0x43, 0x4A, 0x58, 0x22, 0x3B, 0x02, 0x2C, 0x04, 0x23, 0x06,
	0x47, 0x24, 0x36, 0x52, 0x23, 0x1E, 0x10, 0x57, 0x25, 0x75, 0x5F, 0x2D,
	0x0B, 0x5E, 0x74, 0x43, 0x0E, 0x41, 0x40, 0x36, 0x24, 0x51, 0x04, 0x29,
	0x2E, 0x1B, 0x2A, 0x56, 0x1B, 0x1B, 0x1E, 0x37, 0x21, 0x13, 0x32, 0x2E,
	0x25, 0x08, 0x26, 0x34, 0x55, 0x05, 0x38, 0x38, 0x0F, 0x16, 0x08, 0x06,
	0x5D, 0x0B, 0x14, 0x0A, 0x29, 0x2D, 0x04, 0x09, 0x04, 0x2A, 0x00, 0x77,
	0x5A, 0x2B, 0x24, 0x02, 0x1A, 0x26, 0x59, 0x01, 0x01, 0x70, 0x38, 0x07,
	0x59, 0x3A, 0x32, 0x08, 0x0F, 0x17, 0x3F, 0x32, 0x3B, 0x56, 0x25, 0x44,
	0x2D, 0x36, 0x18, 0x22, 0x20, 0x77, 0x24, 0x22, 0x41, 0x19, 0x11, 0x07,
	0x59, 0x25, 0x06, 0x2B, 0x16, 0x20, 0x24, 0x21, 0x73, 0x2A, 0x2F, 0x5B,
	0x33, 0x30, 0x58, 0x24, 0x3B, 0x00, 0x72, 0x2D, 0x10, 0x3D, 0x31, 0x04,
	0x0B, 0x0F, 0x26, 0x12, 0x00, 0x2F, 0x06, 0x04, 0x13, 0x16, 0x2F, 0x2B,
	0x00, 0x04, 0x71, 0x03, 0x0C, 0x2D, 0x3C, 0x11, 0x0F, 0x51, 0x2B, 0x1F,
	0x72, 0x2E, 0x06, 0x2A, 0x32, 0x04, 0x18, 0x2C, 0x5F, 0x31, 0x24, 0x5F,
	0x52, 0x16, 0x19, 0x3B, 0x5B, 0x37, 0x37, 0x52, 0x70, 0x2F, 0x18, 0x19,
	0x38, 0x13, 0x14, 0x03, 0x0F, 0x12, 0x34, 0x00, 0x13, 0x3C, 0x28, 0x05,
	0x59, 0x2F, 0x36, 0x04, 0x0F, 0x27, 0x38, 0x00, 0x1E, 0x34, 0x2F, 0x11,
	0x00, 0x2C, 0x14, 0x19, 0x1B, 0x2A, 0x0F, 0x2A, 0x38, 0x0C, 0x1A, 0x29,
	0x2D, 0x3E, 0x2B, 0x5F, 0x01, 0x05, 0x01, 0x2F, 0x08, 0x24, 0x2A, 0x1C,
	0x56, 0x09, 0x1E, 0x2F, 0x3A, 0x35, 0x39, 0x26, 0x0A, 0x2E, 0x31, 0x0C,
	0x0F, 0x20, 0x05, 0x17, 0x04, 0x28, 0x0B, 0x19, 0x03, 0x5A, 0x21, 0x0C,
	0x3F, 0x00, 0x17, 0x13, 0x1A, 0x3D, 0x2A, 0x3D, 0x13, 0x35, 0x5E, 0x04,
	0x17, 0x02, 0x29, 0x1C, 0x05, 0x2F, 0x25, 0x11, 0x28, 0x2A, 0x2A, 0x0C,
	0x3A, 0x04, 0x30, 0x0C, 0x07, 0x71, 0x5F, 0x2E, 0x5E, 0x12, 0x2A, 0x1C,
	0x19, 0x5A, 0x33, 0x17, 0x07, 0x0F, 0x0C, 0x11, 0x0B, 0x04, 0x31, 0x1E,
	0x0A, 0x3B, 0x1C, 0x02, 0x19, 0x0E, 0x70, 0x24, 0x0A, 0x37, 0x1F, 0x75,
	0x20, 0x3B, 0x41, 0x39, 0x73, 0x54, 0x0A, 0x14, 0x24, 0x0D, 0x5C, 0x30,
	0x06, 0x33, 0x20, 0x15, 0x2F, 0x2D, 0x28, 0x0B, 0x3F, 0x23, 0x36, 0x5A,
	0x38, 0x00, 0x38, 0x3F, 0x26, 0x26, 0x15, 0x00, 0x1A, 0x1D, 0x03, 0x5C,
	0x0F, 0x2A, 0x53, 0x3A, 0x5E, 0x06, 0x09, 0x20, 0x35, 0x20, 0x06, 0x06,
	0x22, 0x2F, 0x3B, 0x38, 0x18, 0x1E, 0x3B, 0x16, 0x18, 0x2F, 0x5F, 0x05,
	0x5B, 0x34, 0x3A, 0x06, 0x38, 0x24, 0x28, 0x41, 0x23, 0x08, 0x1E, 0x0E,
	0x29, 0x28, 0x12, 0x39, 0x0D, 0x26, 0x1D, 0x38, 0x3E, 0x2A, 0x01, 0x05,
	0x76, 0x3A, 0x00, 0x29, 0x3D, 0x2B, 0x5D, 0x51, 0x37, 0x33, 0x29, 0x1E,
	0x58, 0x3D, 0x38, 0x72, 0x38, 0x37, 0x3A, 0x38, 0x30, 0x05, 0x17, 0x1F,
	0x39, 0x75, 0x16, 0x34, 0x58, 0x5E, 0x21, 0x1A, 0x16, 0x34, 0x12, 0x14,
	0x2F, 0x24, 0x16, 0x20, 0x32, 0x24, 0x38, 0x02, 0x09, 0x27, 0x1D, 0x54,
	0x03, 0x04, 0x32, 0x3D, 0x10, 0x58, 0x08, 0x01, 0x14, 0x35, 0x1D, 0x1A,
	0x74, 0x23, 0x14, 0x00, 0x5F, 0x32, 0x00, 0x13, 0x0F, 0x11, 0x6D, 0x2A,
	0x12, 0x5F, 0x58, 0x26, 0x02, 0x12, 0x3B, 0x2A, 0x0D, 0x35, 0x50, 0x03,
	0x32, 0x20, 0x39, 0x28, 0x0F, 0x5A, 0x2F, 0x09, 0x12, 0x18, 0x1E, 0x1A,
	0x2D, 0x11, 0x24, 0x11, 0x76, 0x25, 0x05, 0x2A, 0x3D, 0x36, 0x25, 0x2D,
	0x45, 0x0D, 0x09, 0x5B, 0x25, 0x14, 0x3B, 0x32, 0x2F, 0x13, 0x3E, 0x59,
	0x0C, 0x28, 0x2D, 0x01, 0x02, 0x2E, 0x1E, 0x10, 0x17, 0x11, 0x36, 0x58,
	0x37, 0x01, 0x3B, 0x2E, 0x5F, 0x12, 0x14, 0x1D, 0x35, 0x39, 0x16, 0x58,
	0x23, 0x35, 0x3E, 0x17, 0x34, 0x2A, 0x07, 0x18, 0x0C, 0x5F, 0x3F, 0x0E,
	0x20, 0x23, 0x45, 0x1E, 0x3A, 0x24, 0x2B, 0x41, 0x22, 0x14, 0x2D, 0x29,
	0x0C, 0x5D, 0x08, 0x04, 0x0A, 0x2C, 0x22, 0x29, 0x43, 0x15, 0x28, 0x29,
	0x3A, 0x28, 0x4A, 0x06, 0x09, 0x34, 0x35, 0x29, 0x5F, 0x2F, 0x7B, 0x3D,
	0x07, 0x5A, 0x08, 0x74, 0x3D, 0x27, 0x18, 0x3F, 0x6D, 0x39, 0x12, 0x06,
	0x1E, 0x1B, 0x36, 0x2F, 0x22, 0x23, 0x28, 0x28, 0x08, 0x3C, 0x3C, 0x74,
	0x00, 0x2A, 0x16, 0x27, 0x23, 0x5C, 0x31, 0x57, 0x3E, 0x15, 0x0B, 0x0E,
	0x38, 0x3D, 0x0D, 0x2B, 0x13, 0x0A, 0x1C, 0x24, 0x3A, 0x0E, 0x25, 0x04,
	0x07, 0x2B, 0x23, 0x2B, 0x1A, 0x08, 0x19, 0x10, 0x19, 0x0E, 0x34, 0x19,
	0x17, 0x04, 0x38, 0x73, 0x39, 0x08, 0x2F, 0x00, 0x36, 0x1E, 0x07, 0x2A,
	0x28, 0x75, 0x38, 0x4A, 0x20, 0x0F, 0x6D, 0x03, 0x36, 0x2B, 0x2E, 0x08,
	0x22, 0x08, 0x34, 0x06, 0x06, 0x5D, 0x27, 0x5E, 0x25, 0x06, 0x24, 0x50,
	0x09, 0x33, 0x36, 0x3A, 0x2C, 0x0C, 0x3A, 0x03, 0x39, 0x55, 0x21, 0x53,
	0x17, 0x01, 0x15, 0x25, 0x1B, 0x38, 0x24, 0x55, 0x28, 0x44, 0x33, 0x03,
	0x05, 0x45, 0x0D, 0x7A, 0x3B, 0x2E, 0x24, 0x0C, 0x11, 0x16, 0x20, 0x41,
	0x04, 0x2C, 0x09, 0x28, 0x2C, 0x01, 0x0E, 0x43, 0x39, 0x45, 0x0F, 0x7B,
	0x38, 0x34, 0x05, 0x13, 0x11, 0x39, 0x33, 0x07, 0x5F, 0x14, 0x0A, 0x54,
	0x0A, 0x5A, 0x29, 0x58, 0x59, 0x09, 0x0D, 0x77, 0x3F, 0x18, 0x23, 0x04,
	0x17, 0x27, 0x26, 0x16, 0x03, 0x03, 0x23, 0x54, 0x3B, 0x18, 0x26, 0x2D,
	0x25, 0x3F, 0x03, 0x7A, 0x29, 0x37, 0x59, 0x3E, 0x74, 0x5A, 0x16, 0x2B,
	0x1D, 0x77, 0x24, 0x23, 0x3F, 0x18, 0x15, 0x5A, 0x34, 0x00, 0x39, 0x71,
	0x2F, 0x20, 0x01, 0x29, 0x05, 0x0D, 0x12, 0x1C, 0x0F, 0x14, 0x0F, 0x24,
	0x58, 0x0D, 0x01, 0x3F, 0x12, 0x34, 0x21, 0x01, 0x23, 0x16, 0x16, 0x40,
	0x7B, 0x01, 0x25, 0x37, 0x3A, 0x24, 0x5D, 0x2F, 0x21, 0x04, 0x32, 0x2F,
	0x05, 0x1E, 0x1B, 0x24, 0x06, 0x4E, 0x03, 0x20, 0x7A, 0x19, 0x59, 0x1F,
	0x44, 0x23, 0x0E, 0x59, 0x0D, 0x2D, 0x28, 0x47, 0x30, 0x0C, 0x13, 0x16,
	0x47, 0x37, 0x38, 0x5F, 0x2E, 0x43, 0x2A, 0x18, 0x5F, 0x1A, 0x54, 0x10,
	0x26, 0x59, 0x76, 0x2D, 0x4A, 0x38, 0x58, 0x77, 0x59, 0x2F, 0x2F, 0x24,
	0x12, 0x54, 0x53, 0x3F, 0x3A, 0x74, 0x1F, 0x14, 0x17, 0x38, 0x27, 0x43,
	0x32, 0x05, 0x11, 0x0C, 0x02, 0x06, 0x36, 0x58, 0x1A, 0x5E, 0x2A, 0x02,
	0x1B, 0x69, 0x34, 0x2A, 0x04, 0x21, 0x1B, 0x54, 0x09, 0x5E, 0x25, 0x76,
	0x55, 0x50, 0x08, 0x0C, 0x20, 0x34, 0x23, 0x01, 0x53, 0x24, 0x5C, 0x2B,
	0x23, 0x33, 0x74, 0x28, 0x09, 0x2A, 0x5C, 0x2D, 0x3F, 0x55, 0x28, 0x06,
	0x05, 0x0A, 0x26, 0x02, 0x2A, 0x08, 0x58, 0x10, 0x59, 0x09, 0x13, 0x27,
	0x50, 0x41, 0x5A, 0x38, 0x06, 0x28, 0x3D, 0x5D, 0x20, 0x15, 0x03, 0x5B,
	0x18, 0x17, 0x15, 0x2A, 0x20, 0x1B, 0x2B, 0x26, 0x10, 0x38, 0x18, 0x0A,
	0x0B, 0x04, 0x17, 0x3E, 0x01, 0x0A, 0x58, 0x29, 0x5D, 0x01, 0x09, 0x53,
	0x36, 0x5A, 0x12, 0x34, 0x25, 0x38, 0x27, 0x0F, 0x04, 0x2E, 0x39, 0x1D,
	0x11, 0x1B, 0x4E, 0x27, 0x1E, 0x37, 0x38, 0x4A, 0x3E, 0x40, 0x21, 0x03,
	0x2F, 0x2F, 0x2C, 0x21, 0x05, 0x07, 0x5C, 0x3C, 0x2D, 0x5E, 0x30, 0x39,
	0x22, 0x20, 0x0A, 0x06, 0x57, 0x5C, 0x75, 0x43, 0x54, 0x5C, 0x23, 0x72,
	0x43, 0x59, 0x27, 0x1E, 0x21, 0x21, 0x2D, 0x41, 0x1C, 0x2B, 0x58, 0x16,
	0x06, 0x32, 0x16, 0x0F, 0x03, 0x04, 0x2F, 0x2C, 0x43, 0x19, 0x0C, 0x53,
	0x20, 0x47, 0x32, 0x57, 0x1B, 0x27, 0x27, 0x2C, 0x0C, 0x21, 0x06, 0x58,
	0x30, 0x06, 0x2A, 0x3A, 0x00, 0x2C, 0x2D, 0x40, 0x2A, 0x23, 0x32, 0x2C,
	0x21, 0x36, 0x36, 0x27, 0x56, 0x18, 0x31, 0x1F, 0x3B, 0x1A, 0x1C, 0x25,
	0x54, 0x15, 0x41, 0x3D, 0x11, 0x21, 0x23, 0x2A, 0x21, 0x06, 0x14, 0x31,
	0x19, 0x0C, 0x24, 0x34, 0x22, 0x36, 0x02, 0x04, 0x04, 0x22, 0x0A, 0x21,
	0x37, 0x25, 0x14, 0x2B, 0x1A, 0x72, 0x00, 0x38, 0x3F, 0x08, 0x0B, 0x05,
	0x24, 0x00, 0x21, 0x08, 0x23, 0x28, 0x29, 0x2E, 0x0B, 0x3F, 0x35, 0x5E,
	0x22, 0x33, 0x29, 0x2F, 0x2D, 0x3E, 0x73, 0x26, 0x10, 0x2B, 0x3B, 0x01,
	0x55, 0x06, 0x37, 0x28, 0x34, 0x05, 0x03, 0x06, 0x2A, 0x3A, 0x26, 0x04,
	0x27, 0x0E, 0x04, 0x26, 0x24, 0x1B, 0x5F, 0x2B, 0x58, 0x36, 0x01, 0x38,
	0x14, 0x1C, 0x22, 0x19, 0x02, 0x0B, 0x3E, 0x02, 0x2B, 0x00, 0x76, 0x0B,
	0x38, 0x3F, 0x0C, 0x08, 0x1A, 0x34, 0x06, 0x04, 0x13, 0x5C, 0x2B, 0x3A,
	0x2E, 0x37, 0x1D, 0x30, 0x1D, 0x3B, 0x72, 0x0D, 0x36, 0x3A, 0x5F, 0x08,
	0x24, 0x54, 0x2A, 0x1C, 0x01, 0x0B, 0x0D, 0x3E, 0x00, 0x2C, 0x2D, 0x39,
	0x2D, 0x3D, 0x27, 0x38, 0x12, 0x27, 0x20, 0x07, 0x3E, 0x32, 0x3A, 0x00,
	0x29, 0x02, 0x20, 0x2D, 0x28, 0x17, 0x22, 0x28, 0x58, 0x2E, 0x14, 0x2F,
	0x26, 0x16, 0x20, 0x23, 0x07, 0x0D, 0x2D, 0x23, 0x2A, 0x23, 0x52, 0x5F,
	0x31, 0x12, 0x07, 0x0A, 0x08, 0x2E, 0x06, 0x2F, 0x2A, 0x17, 0x3A, 0x7A,
	0x3F, 0x02, 0x24, 0x0F, 0x08, 0x2A, 0x19, 0x20, 0x1C, 0x25, 0x03, 0x32,
	0x28, 0x1B, 0x05, 0x3D, 0x32, 0x56, 0x22, 0x08, 0x26, 0x20, 0x19, 0x03,
	0x2D, 0x3E, 0x02, 0x24, 0x09, 0x17, 0x04, 0x0E, 0x3D, 0x00, 0x0B, 0x08,
	0x24, 0x1C, 0x31, 0x24, 0x26, 0x02, 0x1D, 0x05, 0x76, 0x3D, 0x2C, 0x3D,
	0x33, 0x2B, 0x24, 0x09, 0x3D, 0x39, 0x0E, 0x19, 0x28, 0x1B, 0x2D, 0x33,
	0x29, 0x0D, 0x0F, 0x3A, 0x31, 0x25, 0x08, 0x2B, 0x33, 0x00, 0x26, 0x2E,
	0x27, 0x2C, 0x07, 0x25, 0x22, 0x0C, 0x5A, 0x0B, 0x0D, 0x24, 0x20, 0x28,
	0x17, 0x14, 0x2D, 0x1F, 0x00, 0x0E, 0x28, 0x58, 0x2D, 0x07, 0x29, 0x47,
	0x22, 0x3C, 0x40, 0x13, 0x54, 0x20, 0x01, 0x21, 0x2B, 0x14, 0x22, 0x41,
	0x0F, 0x32, 0x1B, 0x52, 0x38, 0x09, 0x20, 0x1B, 0x06, 0x28, 0x2F, 0x38,
	0x3C, 0x2E, 0x2B, 0x29, 0x34, 0x1F, 0x56, 0x58, 0x39, 0x29, 0x1A, 0x26,
	0x5F, 0x31, 0x69, 0x08, 0x2F, 0x5A, 0x01, 0x0B, 0x15, 0x2F, 0x45, 0x0E,
	0x13, 0x2F, 0x36, 0x5A, 0x13, 0x17, 0x43, 0x19, 0x05, 0x53, 0x26, 0x06,
	0x4E, 0x45, 0x2C, 0x2C, 0x54, 0x33, 0x45, 0x0E, 0x17, 0x43, 0x58, 0x2A,
	0x0D, 0x2F, 0x07, 0x25, 0x25, 0x3D, 0x71, 0x27, 0x56, 0x08, 0x5E, 0x0E,
	0x5A, 0x31, 0x41, 0x19, 0x77, 0x16, 0x0B, 0x1E, 0x18, 0x25, 0x0A, 0x4E,
	0x45, 0x0D, 0x2C, 0x43, 0x4E, 0x18, 0x5C, 0x24, 0x43, 0x37, 0x1D, 0x5C,
	0x25, 0x5E, 0x06, 0x02, 0x2A, 0x38, 0x26, 0x2C, 0x27, 0x0A, 0x05, 0x0F,
	0x39, 0x58, 0x2A, 0x2A, 0x2D, 0x18, 0x22, 0x2D, 0x2C, 0x5D, 0x13, 0x14,
	0x5C, 0x13, 0x0B, 0x22, 0x2B, 0x04, 0x24, 0x39, 0x2C, 0x2D, 0x12, 0x15,
	0x0B, 0x2F, 0x5B, 0x11, 0x01, 0x38, 0x0B, 0x1C, 0x2F, 0x03, 0x29, 0x0F,
	0x01, 0x1A, 0x6D, 0x03, 0x36, 0x26, 0x2C, 0x32, 0x06, 0x30, 0x45, 0x2E,
	0x7B, 0x0A, 0x11, 0x24, 0x28, 0x08, 0x0E, 0x04, 0x39, 0x04, 0x0B, 0x0B,
	0x54, 0x45, 0x40, 0x6D, 0x25, 0x00, 0x3A, 0x23, 0x30, 0x5D, 0x39, 0x17,
	0x29, 0x14, 0x2F, 0x00, 0x19, 0x58, 0x11, 0x2A, 0x02, 0x3E, 0x58, 0x01,
	0x34, 0x0D, 0x05, 0x2A, 0x27, 0x06, 0x58, 0x0C, 0x0A, 0x20, 0x0F, 0x04,
	0x19, 0x2E, 0x30, 0x38, 0x12, 0x56, 0x08, 0x20, 0x2D, 0x39, 0x3F, 0x0A,
	0x69, 0x2F, 0x0D, 0x2A, 0x12, 0x35, 0x54, 0x13, 0x0C, 0x05, 0x20, 0x22,
	0x31, 0x45, 0x3B, 0x28, 0x04, 0x57, 0x5F, 0x1F, 0x09, 0x03, 0x15, 0x16,
	0x12, 0x34, 0x24, 0x25, 0x58, 0x00, 0x08, 0x3F, 0x12, 0x58, 0x1A, 0x71,
	0x47, 0x53, 0x29, 0x0E, 0x7A, 0x14, 0x2A, 0x0B, 0x01, 0x2C, 0x02, 0x0A,
	0x5B, 0x11, 0x71, 0x02, 0x38, 0x28, 0x5C, 0x24, 0x5F, 0x34, 0x0C, 0x40,
	0x1B, 0x3B, 0x59, 0x0B, 0x25, 0x38, 0x5B, 0x15, 0x20, 0x08, 0x32, 0x43,
	0x4E, 0x1D, 0x5A, 0x25, 0x00, 0x00, 0x1A, 0x1D, 0x2B, 0x43, 0x51, 0x41,
	0x01, 0x71, 0x14, 0x34, 0x1F, 0x59, 0x10, 0x55, 0x51, 0x3E, 0x44, 0x03,
	0x1D, 0x15, 0x18, 0x5E, 0x24, 0x02, 0x0A, 0x18, 0x44, 0x27, 0x0F, 0x11,
	0x39, 0x3A, 0x76, 0x08, 0x2D, 0x25, 0x2E, 0x38, 0x02, 0x22, 0x05, 0x24,
	0x2A, 0x16, 0x4E, 0x1B, 0x01, 0x05, 0x3D, 0x0E, 0x02, 0x09, 0x1B, 0x43,
	0x0F, 0x36, 0x39, 0x20, 0x16, 0x2B, 0x07, 0x06, 0x20, 0x5E, 0x03, 0x59,
	0x32, 0x36, 0x2E, 0x11, 0x3C, 0x19, 0x7B, 0x0E, 0x1B, 0x59, 0x53, 0x73,
	0x5E, 0x52, 0x57, 0x00, 0x34, 0x26, 0x18, 0x14, 0x5A, 0x28, 0x5F, 0x36,
	0x17, 0x12, 0x30, 0x2D, 0x07, 0x27, 0x44, 0x23, 0x1E, 0x25, 0x08, 0x07,
	0x7A, 0x3D, 0x24, 0x57, 0x1E, 0x26, 0x3F, 0x25, 0x2C, 0x5D, 0x31, 0x3B,
	0x23, 0x25, 0x12, 0x7A, 0x29, 0x2F, 0x2A, 0x44, 0x3B, 0x0D, 0x00, 0x58,
	0x2A, 0x07, 0x1C, 0x23, 0x5E, 0x53, 0x31, 0x3A, 0x58, 0x0B, 0x5B, 0x00,
	0x5C, 0x55, 0x20, 0x19, 0x69, 0x3B, 0x19, 0x08, 0x13, 0x7A, 0x2D, 0x0F,
	0x57, 0x3B, 0x3B, 0x1E, 0x39, 0x41, 0x33, 0x16, 0x2D, 0x0F, 0x1B, 0x05,
	0x3A, 0x43, 0x09, 0x38, 0x52, 0x14, 0x1B, 0x05, 0x1B, 0x23, 0x26, 0x08,
	0x0B, 0x56, 0x23, 0x1A, 0x1E, 0x1B, 0x3F, 0x2E, 0x7B, 0x04, 0x53, 0x5B,
	0x53, 0x37, 0x3C, 0x2C, 0x58, 0x0A, 0x30, 0x21, 0x0B, 0x36, 0x2D, 0x2C,
	0x5F, 0x0D, 0x05, 0x07, 0x27, 0x38, 0x2B, 0x08, 0x06, 0x12, 0x3E, 0x18,
	0x41, 0x3F, 0x23, 0x09, 0x1B, 0x5C, 0x38, 0x34, 0x0E, 0x35, 0x58, 0x09,
	0x7B, 0x5E, 0x0A, 0x3A, 0x26, 0x75, 0x43, 0x2E, 0x45, 0x23, 0x12, 0x06,
	0x17, 0x00, 0x1F, 0x0F, 0x3A, 0x14, 0x26, 0x3D, 0x70, 0x3C, 0x2F, 0x18,
	0x52, 0x0B, 0x26, 0x36, 0x16, 0x44, 0x2F, 0x55, 0x31, 0x34, 0x1C, 0x10,
	0x29, 0x29, 0x3A, 0x0E, 0x0F, 0x0A, 0x2D, 0x38, 0x39, 0x32, 0x3B, 0x22,
	0x01, 0x27, 0x2B, 0x5D, 0x23, 0x41, 0x32, 0x12, 0x27, 0x15, 0x5E, 0x09,
	0x08, 0x27, 0x09, 0x0C, 0x1F, 0x7B, 0x0E, 0x4A, 0x5C, 0x09, 0x0D, 0x0B,
	0x14, 0x3C, 0x5F, 0x1A, 0x5D, 0x38, 0x01, 0x06, 0x7B, 0x2E, 0x57, 0x5B,
	0x3B, 0x0E, 0x02, 0x0E, 0x00, 0x2E, 0x75, 0x1A, 0x51, 0x3D, 0x25, 0x12,
	0x43, 0x56, 0x17, 0x0D, 0x72, 0x54, 0x20, 0x1B, 0x2C, 0x70, 0x00, 0x39,
	0x1B, 0x26, 0x25, 0x1B, 0x59, 0x21, 0x01, 0x10, 0x07, 0x37, 0x59, 0x08,
	0x69, 0x59, 0x0C, 0x34, 0x29, 0x7B, 0x5A, 0x2E, 0x18, 0x23, 0x0E, 0x2E,
	0x02, 0x20, 0x09, 0x0F, 0x3E, 0x4A, 0x0F, 0x01, 0x24, 0x24, 0x57, 0x37,
	0x3F, 0x05, 0x1B, 0x19, 0x29, 0x3F, 0x36, 0x1D, 0x10, 0x5C, 0x0D, 0x1B,
	0x35, 0x4E, 0x1B, 0x1C, 0x3B, 0x00, 0x24, 0x29, 0x1C, 0x17, 0x43, 0x29,
	0x0B, 0x02, 0x15, 0x0A, 0x29, 0x3C, 0x3C, 0x16, 0x1F, 0x2E, 0x1E, 0x0F,
	0x21, 0x23, 0x29, 0x36, 0x3E, 0x14, 0x00, 0x37, 0x17, 0x1F, 0x3A, 0x5D,
	0x58, 0x5C, 0x13, 0x18, 0x43, 0x09, 0x57, 0x1A, 0x2C, 0x06, 0x54, 0x1A,
	0x38, 0x15, 0x25, 0x3B, 0x59, 0x0D, 0x2C, 0x3D, 0x05, 0x56, 0x27, 0x16,
	0x1C, 0x00, 0x14, 0x0E, 0x09, 0x5B, 0x2C, 0x5D, 0x02, 0x34, 0x1C, 0x04,
	0x34, 0x08, 0x73, 0x06, 0x11, 0x56, 0x13, 0x0F, 0x59, 0x50, 0x21, 0x28,
	0x12, 0x5F, 0x51, 0x0A, 0x5B, 0x17, 0x25, 0x2B, 0x0A, 0x3A, 0x34, 0x01,
	0x15, 0x56, 0x5A, 0x7B, 0x0F, 0x0B, 0x0F, 0x39, 0x05, 0x14, 0x1B, 0x5A,
	0x58, 0x14, 0x5F, 0x0F, 0x5C, 0x26, 0x6D, 0x5D, 0x16, 0x3D, 0x0A, 0x16,
	0x5A, 0x57, 0x5B, 0x31, 0x2C, 0x0E, 0x06, 0x38, 0x1D, 0x05, 0x0D, 0x11,
	0x3C, 0x5F, 0x00, 0x1B, 0x09, 0x5D, 0x31, 0x0B, 0x54, 0x11, 0x1F, 0x05,
	0x70, 0x47, 0x12, 0x05, 0x1D, 0x2B, 0x2B, 0x04, 0x1A, 0x0D, 0x21, 0x0E,
	0x0B, 0x57, 0x19, 0x29, 0x04, 0x0C, 0x07, 0x5E, 0x0E, 0x59, 0x10, 0x3A,
	0x44, 0x2F, 0x5D, 0x29, 0x17, 0x2C, 0x23, 0x43, 0x4A, 0x5F, 0x40, 0x2F,
	0x55, 0x39, 0x05, 0x08, 0x0F, 0x01, 0x4E, 0x06, 0x2F, 0x26, 0x24, 0x57,
	0x2A, 0x3F, 0x73, 0x2F, 0x25, 0x16, 0x5F, 0x08, 0x21, 0x11, 0x2D, 0x1C,
	0x15, 0x27, 0x27, 0x58, 0x03, 0x28, 0x1D, 0x17, 0x29, 0x05, 0x26, 0x3C,
	0x22, 0x45, 0x59, 0x3A, 0x38, 0x26, 0x41, 0x11, 0x77, 0x08, 0x57, 0x26,
	0x3A, 0x31, 0x0A, 0x2B, 0x0C, 0x1F, 0x23, 0x0A, 0x36, 0x1A, 0x53, 0x23,
	0x19, 0x14, 0x16, 0x3E, 0x70, 0x09, 0x31, 0x2A, 0x01, 0x0A, 0x59, 0x09,
	0x3B, 0x59, 0x72, 0x24, 0x52, 0x0C, 0x3D, 0x1B, 0x29, 0x09, 0x3B, 0x3C,
	0x6D, 0x43, 0x52, 0x1A, 0x5D, 0x06, 0x0F, 0x4E, 0x34, 0x04, 0x24, 0x5D,
	0x39, 0x1B, 0x3C, 0x3B, 0x1B, 0x2E, 0x04, 0x29, 0x74, 0x0E, 0x23, 0x2B,
	0x0D, 0x69, 0x3B, 0x53, 0x5B, 0x3E, 0x23, 0x0A, 0x16, 0x1F, 0x31, 0x07,
	0x39, 0x30, 0x41, 0x03, 0x76, 0x1B, 0x00, 0x3E, 0x11, 0x2D, 0x03, 0x57,
	0x01, 0x44, 0x21, 0x03, 0x2D, 0x5C, 0x2D, 0x72, 0x5F, 0x36, 0x2D, 0x05,
	0x23, 0x26, 0x2C, 0x02, 0x28, 0x72, 0x08, 0x31, 0x0A, 0x1A, 0x75, 0x09,
	0x4E, 0x18, 0x2F, 0x76, 0x04, 0x05, 0x29, 0x31, 0x73, 0x3B, 0x2C, 0x1B,
	0x0A, 0x24, 0x0E, 0x20, 0x19, 0x06, 0x34, 0x0A, 0x53, 0x34, 0x12, 0x31,
	0x5A, 0x2E, 0x5E, 0x3E, 0x75, 0x1E, 0x56, 0x1C, 0x0A, 0x00, 0x0D, 0x4E,
	0x08, 0x58, 0x32, 0x58, 0x03, 0x0F, 0x12, 0x14, 0x23, 0x08, 0x5F, 0x01,
	0x16, 0x34, 0x0B, 0x08, 0x1B, 0x2B, 0x23, 0x02, 0x02, 0x1D, 0x1A, 0x34,
	0x16, 0x56, 0x5A, 0x06, 0x20, 0x24, 0x57, 0x1F, 0x29, 0x27, 0x09, 0x28,
	0x5C, 0x05, 0x3F, 0x4E, 0x5D, 0x11, 0x14, 0x02, 0x0D, 0x5F, 0x0E, 0x07,
	0x3A, 0x0C, 0x26, 0x26, 0x12, 0x16, 0x53, 0x1A, 0x29, 0x10, 0x2B, 0x09,
	0x0D, 0x3F, 0x37, 0x00, 0x55, 0x57, 0x18, 0x70, 0x3E, 0x18, 0x3A, 0x1F,
	0x20, 0x5C, 0x0E, 0x3B, 0x0D, 0x20, 0x58, 0x07, 0x37, 0x31, 0x32, 0x08,
	0x2E, 0x5F, 0x5C, 0x7B, 0x1D, 0x29, 0x58, 0x00, 0x00, 0x0F, 0x17, 0x57,
	0x04, 0x01, 0x3D, 0x15, 0x23, 0x25, 0x08, 0x01, 0x1B, 0x0D, 0x11, 0x73,
	0x19, 0x52, 0x19, 0x27, 0x0B, 0x1B, 0x17, 0x3E, 0x27, 0x0E, 0x38, 0x38,
	0x29, 0x09, 0x13, 0x1A, 0x2C, 0x1B, 0x5C, 0x28, 0x3A, 0x57, 0x59, 0x13,
	0x34, 0x09, 0x04, 0x3C, 0x0C, 0x29, 0x00, 0x37, 0x1D, 0x5B, 0x72, 0x34,
	0x58, 0x27, 0x06, 0x11, 0x2E, 0x14, 0x14, 0x1D, 0x7A, 0x09, 0x29, 0x1B,
	0x5D, 0x09, 0x06, 0x50, 0x16, 0x0C, 0x2C, 0x5F, 0x52, 0x01, 0x3F, 0x12,
	0x05, 0x2D, 0x1E, 0x04, 0x2F, 0x02, 0x05, 0x57, 0x40, 0x76, 0x18, 0x0B,
	0x3B, 0x38, 0x0F, 0x21, 0x09, 0x07, 0x39, 0x24, 0x15, 0x0F, 0x5A, 0x33,
	0x32, 0x08, 0x31, 0x05, 0x5C, 0x0C, 0x00, 0x4A, 0x5C, 0x38, 0x08, 0x0D,
	0x31, 0x58, 0x3F, 0x29, 0x1F, 0x10, 0x08, 0x58, 0x37, 0x23, 0x09, 0x22,
	0x1E, 0x25, 0x5D, 0x13, 0x2C, 0x1A, 0x30, 0x22, 0x08, 0x5C, 0x5E, 0x24,
	0x09, 0x25, 0x59, 0x3A, 0x20, 0x19, 0x32, 0x5B, 0x0A, 0x07, 0x47, 0x31,
	0x1F, 0x1F, 0x28, 0x06, 0x2A, 0x59, 0x52, 0x04, 0x1C, 0x54, 0x09, 0x09,
	0x14, 0x24, 0x50, 0x0F, 0x31, 0x3A, 0x08, 0x35, 0x41, 0x2E, 0x6D, 0x3C,
	0x06, 0x37, 0x20, 0x0E, 0x15, 0x35, 0x26, 0x25, 0x72, 0x00, 0x37, 0x18,
	0x0A, 0x06, 0x47, 0x39, 0x16, 0x08, 0x38, 0x36, 0x36, 0x41, 0x3B, 0x08,
	0x15, 0x10, 0x1D, 0x40, 0x77, 0x1F, 0x50, 0x5A, 0x39, 0x7A, 0x2B, 0x23,
	0x37, 0x24, 0x17, 0x14, 0x26, 0x0D, 0x5E, 0x1B, 0x36, 0x35, 0x45, 0x59,
	0x69, 0x59, 0x09, 0x14, 0x1D, 0x36, 0x06, 0x29, 0x57, 0x28, 0x0D, 0x54,
	0x2C, 0x0D, 0x0E, 0x31, 0x05, 0x15, 0x5E, 0x0E, 0x1A, 0x55, 0x59, 0x19,
	0x31, 0x30, 0x28, 0x35, 0x5C, 0x1D, 0x0C, 0x5F, 0x57, 0x1E, 0x19, 0x05,
	0x23, 0x31, 0x1D, 0x1C, 0x7A, 0x43, 0x32, 0x45, 0x5D, 0x7A, 0x3E, 0x36,
	0x39, 0x5A, 0x33, 0x5F, 0x17, 0x01, 0x11, 0x38, 0x05, 0x52, 0x5D, 0x23,
	0x20, 0x55, 0x15, 0x01, 0x5F, 0x18, 0x3D, 0x39, 0x1B, 0x58, 0x0C, 0x19,
	0x25, 0x1D, 0x58, 0x15, 0x36, 0x50, 0x08, 0x18, 0x18, 0x36, 0x2F, 0x1A,
	0x5D, 0x11, 0x09, 0x0A, 0x04, 0x59, 0x0C, 0x24, 0x13, 0x2A, 0x3E, 0x7A,
	0x47, 0x53, 0x1E, 0x52, 0x38, 0x5B, 0x26, 0x06, 0x0F, 0x11, 0x0D, 0x07,
	0x20, 0x00, 0x37, 0x2F, 0x19, 0x14, 0x19, 0x72, 0x18, 0x07, 0x18, 0x20,
	0x38, 0x26, 0x51, 0x45, 0x1F, 0x31, 0x05, 0x59, 0x19, 0x27, 0x15, 0x5F,
	0x51, 0x0B, 0x2C, 0x3A, 0x1D, 0x57, 0x5D, 0x23, 0x17, 0x3E, 0x31, 0x18,
	0x1D, 0x00, 0x03, 0x56, 0x41, 0x08, 0x21, 0x35, 0x17, 0x5E, 0x20, 0x73,
	0x43, 0x14, 0x23, 0x59, 0x06, 0x20, 0x2F, 0x0A, 0x1E, 0x0A, 0x26, 0x53,
	0x57, 0x27, 0x25, 0x59, 0x26, 0x1D, 0x24, 0x0D, 0x47, 0x27, 0x00, 0x3B,
	0x05, 0x0E, 0x07, 0x05, 0x40, 0x26, 0x01, 0x28, 0x05, 0x38, 0x37, 0x1E,
	0x19, 0x5D, 0x05, 0x11, 0x28, 0x51, 0x00, 0x01, 0x09, 0x26, 0x4E, 0x26,
	0x29, 0x15, 0x55, 0x54, 0x5E, 0x1F, 0x69, 0x1C, 0x05, 0x2B, 0x02, 0x21,
	0x34, 0x05, 0x2D, 0x3D, 0x10, 0x3B, 0x12, 0x0A, 0x59, 0x0A, 0x29, 0x27,
	0x0A, 0x58, 0x70, 0x23, 0x2C, 0x0F, 0x08, 0x37, 0x05, 0x09, 0x1D, 0x33,
	0x30, 0x1A, 0x4A, 0x17, 0x5A, 0x7A, 0x23, 0x2D, 0x0D, 0x0D, 0x2F, 0x2F,
	0x34, 0x3F, 0x58, 0x18, 0x00, 0x56, 0x2A, 0x13, 0x0F, 0x3B, 0x24, 0x3E,
	0x3D, 0x0B, 0x20, 0x03, 0x00, 0x08, 0x18, 0x02, 0x31, 0x38, 0x58, 0x07,
	0x0E, 0x31, 0x0F, 0x08, 0x0D, 0x3C, 0x56, 0x1D, 0x19, 0x34, 0x24, 0x36,
	0x21, 0x5A, 0x0E, 0x3B, 0x0B, 0x06, 0x0D, 0x73, 0x23, 0x14, 0x09, 0x3C,
	0x17, 0x5F, 0x19, 0x04, 0x1D, 0x06, 0x5B, 0x56, 0x1D, 0x3E, 0x30, 0x3B,
	0x36, 0x18, 0x3E, 0x08, 0x5E, 0x16, 0x1B, 0x28, 0x38, 0x0A, 0x53, 0x38,
	0x1D, 0x11, 0x0F, 0x51, 0x5D, 0x00, 0x70, 0x1B, 0x0B, 0x1F, 0x22, 0x09,
	0x26, 0x50, 0x14, 0x3C, 0x12, 0x59, 0x2A, 0x5D, 0x3F, 0x15, 0x34, 0x13,
	0x06, 0x20, 0x29, 0x14, 0x2D, 0x5D, 0x1B, 0x07, 0x21, 0x33, 0x57, 0x24,
	0x70, 0x20, 0x51, 0x5A, 0x11, 0x0F, 0x0D, 0x54, 0x5D, 0x28, 0x00, 0x47,
	0x52, 0x3E, 0x2C, 0x2C, 0x47, 0x05, 0x21, 0x11, 0x2F, 0x0A, 0x29, 0x56,
	0x5A, 0x34, 0x24, 0x26, 0x29, 0x40, 0x1B, 0x39, 0x19, 0x3F, 0x44, 0x23,
	0x5B, 0x4E, 0x26, 0x06, 0x15, 0x0F, 0x4E, 0x57, 0x53, 0x27, 0x43, 0x08,
	0x5F, 0x3F, 0x0F, 0x09, 0x52, 0x00, 0x53, 0x10, 0x43, 0x59, 0x41, 0x03,
	0x11, 0x58, 0x18, 0x37, 0x06, 0x71, 0x5C, 0x35, 0x3E, 0x04, 0x23, 0x1A,
	0x0A, 0x3B, 0x39, 0x34, 0x28, 0x24, 0x41, 0x32, 0x0D, 0x5E, 0x08, 0x03,
	0x11, 0x1B, 0x5A, 0x30, 0x03, 0x0A, 0x00, 0x5F, 0x36, 0x26, 0x19, 0x07,
	0x55, 0x25, 0x45, 0x39, 0x2D, 0x20, 0x30, 0x05, 0x1F, 0x28, 0x38, 0x29,
	0x45, 0x33, 0x71, 0x2F, 0x0C, 0x3C, 0x53, 0x7A, 0x05, 0x19, 0x1D, 0x5A,
	0x03, 0x55, 0x0A, 0x08, 0x1D, 0x73, 0x47, 0x18, 0x2B, 0x3A, 0x34, 0x05,
	0x53, 0x26, 0x06, 0x04, 0x25, 0x51, 0x5A, 0x5F, 0x73, 0x54, 0x50, 0x04,
	0x25, 0x7A, 0x0E, 0x2F, 0x26, 0x0E, 0x30, 0x02, 0x02, 0x34, 0x5D, 0x36,
	0x59, 0x03, 0x3A, 0x44, 0x3B, 0x43, 0x36, 0x58, 0x5C, 0x69, 0x15, 0x3B,
	0x39, 0x3B, 0x71, 0x07, 0x51, 0x18, 0x23, 0x70, 0x05, 0x37, 0x1B, 0x13,
	0x72, 0x01, 0x39, 0x3E, 0x2F, 0x2C, 0x2D, 0x32, 0x0C, 0x59, 0x06, 0x3C,
	0x3B, 0x25, 0x09, 0x7B, 0x3A, 0x18, 0x3D, 0x3C, 0x72, 0x18, 0x4E, 0x2B,
	0x39, 0x71, 0x15, 0x10, 0x3A, 0x52, 0x35, 0x03, 0x07, 0x0B, 0x06, 0x74,
	0x14, 0x38, 0x29, 0x0A, 0x26, 0x24, 0x39, 0x57, 0x26, 0x72, 0x0E, 0x55,
	0x38, 0x22, 0x69, 0x07, 0x57, 0x1C, 0x27, 0x26, 0x2B, 0x30, 0x18, 0x06,
	0x18, 0x05, 0x02, 0x5B, 0x1B, 0x09, 0x58, 0x28, 0x17, 0x25, 0x34, 0x43,
	0x37, 0x5F, 0x20, 0x75, 0x18, 0x4A, 0x45, 0x32, 0x74, 0x23, 0x03, 0x0C,
	0x38, 0x15, 0x1A, 0x32, 0x1C, 0x27, 0x76, 0x58, 0x25, 0x57, 0x3D, 0x0C,
	0x3C, 0x0D, 0x41, 0x11, 0x13, 0x09, 0x0B, 0x00, 0x5D, 0x32, 0x47, 0x02,
	0x1A, 0x52, 0x7A, 0x19, 0x52, 0x24, 0x28, 0x10, 0x02, 0x19, 0x14, 0x0F,
	0x24, 0x28, 0x16, 0x02, 0x0F, 0x34, 0x24, 0x14, 0x34, 0x29, 0x21, 0x18,
	0x0D, 0x45, 0x32, 0x34, 0x26, 0x54, 0x5A, 0x00, 0x69, 0x54, 0x52, 0x5F,
	0x0A, 0x3A, 0x20, 0x15, 0x20, 0x24, 0x1B, 0x35, 0x22, 0x07, 0x21, 0x06,
	0x1E, 0x0B, 0x0B, 0x2D, 0x21, 0x2A, 0x56, 0x38, 0x0D, 0x36, 0x3D, 0x15,
	0x2A, 0x38, 0x38, 0x04, 0x32, 0x22, 0x44, 0x23, 0x2B, 0x52, 0x28, 0x26,
	0x33, 0x06, 0x0B, 0x1D, 0x1D, 0x09, 0x27, 0x19, 0x24, 0x53, 0x73, 0x09,
	0x02, 0x14, 0x1C, 0x73, 0x59, 0x56, 0x37, 0x5A, 0x1A, 0x19, 0x4A, 0x08,
	0x04, 0x2C, 0x3A, 0x0D, 0x5D, 0x5D, 0x0A, 0x20, 0x12, 0x5C, 0x21, 0x11,
	0x59, 0x0A, 0x58, 0x27, 0x24, 0x15, 0x10, 0x0C, 0x3C, 0x08, 0x5B, 0x18,
	0x0A, 0x08, 0x69, 0x14, 0x50, 0x19, 0x53, 0x16, 0x0D, 0x50, 0x22, 0x08,
	0x14, 0x07, 0x50, 0x56, 0x1E, 0x27, 0x38, 0x56, 0x5B, 0x5E, 0x13, 0x36,
	0x4E, 0x1A, 0x39, 0x2C, 0x04, 0x34, 0x0B, 0x23, 0x32, 0x18, 0x55, 0x37,
	0x24, 0x15, 0x2E, 0x52, 0x16, 0x3E, 0x26, 0x5E, 0x10, 0x1C, 0x01, 0x34,
	0x1D, 0x56, 0x26, 0x5C, 0x08, 0x05, 0x50, 0x21, 0x09, 0x16, 0x34, 0x07,
	0x41, 0x26, 0x77, 0x39, 0x54, 0x5D, 0x20, 0x33, 0x3D, 0x00, 0x5B, 0x0A,
	0x38, 0x3C, 0x37, 0x34, 0x0E, 0x0C, 0x1D, 0x15, 0x06, 0x39, 0x27, 0x24,
	0x10, 0x1C, 0x3E, 0x74, 0x1C, 0x53, 0x02, 0x5C, 0x6D, 0x24, 0x32, 0x57,
	0x12, 0x0F, 0x00, 0x28, 0x37, 0x44, 0x33, 0x5F, 0x2B, 0x58, 0x5F, 0x70,
	0x3B, 0x54, 0x0D, 0x59, 0x7B, 0x19, 0x00, 0x24, 0x5C, 0x70, 0x3B, 0x11,
	0x20, 0x52, 0x12, 0x5E, 0x0B, 0x1A, 0x1C, 0x77, 0x23, 0x03, 0x38, 0x0A,
	0x0B, 0x5F, 0x50, 0x5D, 0x12, 0x0B, 0x58, 0x05, 0x14, 0x3D, 0x1A, 0x09,
	0x57, 0x39, 0x26, 0x16, 0x0E, 0x58, 0x5E, 0x12, 0x24, 0x05, 0x27, 0x23,
	0x0D, 0x69, 0x0A, 0x19, 0x1A, 0x44, 0x18, 0x28, 0x4A, 0x1C, 0x09, 0x72,
	0x3E, 0x17, 0x45, 0x5A, 0x23, 0x36, 0x2D, 0x27, 0x5E, 0x2C, 0x3F, 0x15,
	0x58, 0x2F, 0x30, 0x0A, 0x39, 0x0B, 0x06, 0x05, 0x29, 0x4A, 0x0A, 0x06,
	0x16, 0x20, 0x54, 0x1B, 0x3E, 0x2A, 0x03, 0x51, 0x3B, 0x0A, 0x03, 0x3F,
	0x18, 0x58, 0x3A, 0x6D, 0x01, 0x1B, 0x1E, 0x39, 0x75, 0x3F, 0x58, 0x36,
	0x0A, 0x74, 0x0F, 0x52, 0x45, 0x12, 0x26, 0x1D, 0x0D, 0x24, 0x0E, 0x77,
	0x58, 0x00, 0x5D, 0x38, 0x2B, 0x0D, 0x18, 0x5D, 0x06, 0x70, 0x36, 0x34,
	0x39, 0x5E, 0x2A, 0x00, 0x53, 0x2B, 0x3D, 0x20, 0x0A, 0x0D, 0x17, 0x0A,
	0x05, 0x59, 0x27, 0x16, 0x27, 0x0F, 0x3C, 0x23, 0x08, 0x06, 0x30, 0x39,
	0x13, 0x27, 0x13, 0x36, 0x27, 0x0D, 0x20, 0x44, 0x12, 0x1C, 0x09, 0x5A,
	0x26, 0x2F, 0x22, 0x16, 0x23, 0x06, 0x6D, 0x2F, 0x2B, 0x0F, 0x3E, 0x12,
	0x2B, 0x02, 0x58, 0x0E, 0x2F, 0x05, 0x54, 0x28, 0x31, 0x35, 0x36, 0x0D,
	0x3A, 0x1F, 0x27, 0x1D, 0x2E, 0x2A, 0x3B, 0x69, 0x1B, 0x31, 0x04, 0x26,
	0x23, 0x5B, 0x37, 0x1B, 0x12, 0x76, 0x55, 0x36, 0x14, 0x18, 0x7A, 0x54,
	0x4E, 0x41, 0x3C, 0x7A, 0x08, 0x55, 0x1A, 0x3F, 0x20, 0x0D, 0x3B, 0x1C,
	0x3D, 0x14, 0x1A, 0x0D, 0x2F, 0x20, 0x15, 0x0A, 0x0C, 0x3F, 0x26, 0x07,
	0x27, 0x1B, 0x17, 0x02, 0x69, 0x16, 0x0D, 0x05, 0x1F, 0x1B, 0x0E, 0x57,
	0x36, 0x1F, 0x2B, 0x47, 0x2F, 0x3D, 0x33, 0x30, 0x47, 0x3B, 0x3E, 0x5E,
	0x3A, 0x5F, 0x11, 0x2B, 0x19, 0x31, 0x16, 0x2A, 0x18, 0x01, 0x0E, 0x21,
	0x14, 0x0B, 0x27, 0x03, 0x18, 0x32, 0x17, 0x1F, 0x2F, 0x18, 0x0A, 0x5F,
	0x0E, 0x6D, 0x19, 0x11, 0x0D, 0x24, 0x24, 0x15, 0x13, 0x3C, 0x5A, 0x0C,
	0x18, 0x16, 0x5D, 0x01, 0x0E, 0x07, 0x17, 0x57, 0x53, 0x16, 0x2E, 0x59,
	0x5B, 0x28, 0x16, 0x19, 0x50, 0x29, 0x05, 0x24, 0x00, 0x56, 0x16, 0x32,
	0x37, 0x36, 0x29, 0x59, 0x00, 0x12, 0x5E, 0x15, 0x1D, 0x21, 0x6D, 0x15,
	0x39, 0x0B, 0x5C, 0x13, 0x1B, 0x14, 0x21, 0x1D, 0x04, 0x16, 0x56, 0x39,
	0x5E, 0x27, 0x3B, 0x12, 0x14, 0x29, 0x28, 0x1F, 0x51, 0x34, 0x1D, 0x00,
	0x3B, 0x50, 0x07, 0x02, 0x21, 0x00, 0x20, 0x1A, 0x08, 0x16, 0x20, 0x31,
	0x3B, 0x52, 0x7B, 0x54, 0x24, 0x1F, 0x25, 0x35, 0x28, 0x4A, 0x57, 0x12,
	0x28, 0x5A, 0x18, 0x41, 0x2D, 0x74, 0x55, 0x59, 0x17, 0x1B, 0x31, 0x0D,
	0x37, 0x5F, 0x0F, 0x7A, 0x43, 0x28, 0x16, 0x21, 0x7B, 0x00, 0x39, 0x5D,
	0x1C, 0x34, 0x1D, 0x0E, 0x36, 0x06, 0x0A, 0x36, 0x07, 0x1C, 0x25, 0x15,
	0x47, 0x13, 0x08, 0x38, 0x11, 0x5B, 0x2C, 0x04, 0x1F, 0x77, 0x5C, 0x19,
	0x29, 0x06, 0x2A, 0x5D, 0x2B, 0x22, 0x1F, 0x2E, 0x03, 0x05, 0x23, 0x20,
	0x2C, 0x19, 0x23, 0x20, 0x1F, 0x36, 0x59, 0x58, 0x1C, 0x25, 0x32, 0x05,
	0x18, 0x5A, 0x29, 0x08, 0x5C, 0x38, 0x37, 0x40, 0x7B, 0x1E, 0x03, 0x14,
	0x13, 0x72, 0x16, 0x2A, 0x07, 0x21, 0x71, 0x5F, 0x59, 0x45, 0x02, 0x2A,
	0x05, 0x0A, 0x02, 0x3B, 0x20, 0x07, 0x50, 0x45, 0x5F, 0x0D, 0x3E, 0x16,
	0x34, 0x1F, 0x09, 0x55, 0x02, 0x1E, 0x26, 0x27, 0x22, 0x04, 0x5F, 0x0D,
	0x08, 0x07, 0x36, 0x56, 0x3C, 0x75, 0x23, 0x22, 0x5D, 0x59, 0x75, 0x22,
	0x17, 0x41, 0x23, 0x18, 0x0E, 0x54, 0x5D, 0x1A, 0x33, 0x39, 0x32, 0x45,
	0x40, 0x0D, 0x22, 0x22, 0x56, 0x3A, 0x1A, 0x19, 0x24, 0x18, 0x5E, 0x70,
	0x47, 0x53, 0x45, 0x1F, 0x17, 0x5C, 0x03, 0x45, 0x11, 0x26, 0x09, 0x2C,
	0x22, 0x13, 0x01, 0x39, 0x09, 0x17, 0x0C, 0x08, 0x43, 0x12, 0x5A, 0x31,
	0x14, 0x5E, 0x4E, 0x5D, 0x59, 0x07, 0x39, 0x16, 0x22, 0x31, 0x09, 0x1A,
	0x07, 0x29, 0x21, 0x77, 0x1C, 0x10, 0x2C, 0x0E, 0x15, 0x22, 0x17, 0x41,
	0x3E, 0x12, 0x21, 0x57, 0x09, 0x33, 0x08, 0x58, 0x4E, 0x18, 0x32, 0x2C,
	0x35, 0x19, 0x01, 0x2D, 0x0F, 0x16, 0x03, 0x28, 0x27, 0x0D, 0x5B, 0x1B,
	0x3C, 0x07, 0x0C, 0x03, 0x36, 0x3E, 0x0D, 0x77, 0x43, 0x08, 0x3D, 0x39,
	0x28, 0x55, 0x23, 0x5A, 0x18, 0x28, 0x28, 0x10, 0x3D, 0x04, 0x0C, 0x25,
	0x14, 0x26, 0x19, 0x32, 0x18, 0x3B, 0x08, 0x3F, 0x03, 0x1E, 0x02, 0x22,
	0x00, 0x70, 0x3D, 0x50, 0x2A, 0x05, 0x37, 0x5D, 0x29, 0x09, 0x06, 0x0A,
	0x02, 0x19, 0x24, 0x26, 0x34, 0x3E, 0x58, 0x1F, 0x21, 0x0C, 0x20, 0x02,
	0x26, 0x0D, 0x20, 0x1B, 0x19, 0x01, 0x0A, 0x10, 0x03, 0x15, 0x3D, 0x18,
	0x69, 0x36, 0x10, 0x0D, 0x3F, 0x21, 0x3B, 0x08, 0x5E, 0x59, 0x33, 0x59,
	0x28, 0x0B, 0x5A, 0x1A, 0x28, 0x55, 0x04, 0x0E, 0x1A, 0x38, 0x33, 0x56,
	0x44, 0x08, 0x3C, 0x18, 0x3B, 0x1F, 0x16, 0x35, 0x1B, 0x1A, 0x1B, 0x18,
	0x59, 0x24, 0x18, 0x3B, 0x2F, 0x09, 0x2E, 0x5F, 0x0F, 0x2D, 0x14, 0x11,
	0x3C, 0x2C, 0x11, 0x23, 0x03, 0x3B, 0x01, 0x26, 0x5A, 0x53, 0x0B, 0x1B,
	0x76, 0x1C, 0x19, 0x04, 0x5C, 0x0F, 0x07, 0x35, 0x26, 0x5A, 0x23, 0x0A,
	0x18, 0x04, 0x2E, 0x33, 0x02, 0x2D, 0x20, 0x40, 0x3B, 0x23, 0x51, 0x3E,
	0x24, 0x15, 0x22, 0x39, 0x5C, 0x00, 0x32, 0x15, 0x13, 0x02, 0x19, 0x2F,
	0x36, 0x11, 0x0A, 0x53, 0x36, 0x58, 0x57, 0x05, 0x13, 0x0D, 0x0F, 0x2E,
	0x0A, 0x2F, 0x2B, 0x14, 0x51, 0x04, 0x29, 0x3A, 0x3D, 0x04, 0x58, 0x0E,
	0x2D, 0x00, 0x05, 0x00, 0x07, 0x2C, 0x02, 0x34, 0x5B, 0x08, 0x23, 0x18,
	0x07, 0x1B, 0x23, 0x29, 0x24, 0x05, 0x3D, 0x0E, 0x69, 0x5B, 0x37, 0x29,
	0x1F, 0x73, 0x43, 0x05, 0x3E, 0x1C, 0x77, 0x59, 0x37, 0x3C, 0x53, 0x2B,
	0x1E, 0x35, 0x17, 0x59, 0x32, 0x19, 0x3B, 0x1A, 0x1F, 0x0C, 0x19, 0x53,
	0x08, 0x52, 0x23, 0x2F, 0x37, 0x36, 0x06, 0x32, 0x29, 0x51, 0x34, 0x06,
	0x0D, 0x14, 0x02, 0x5E, 0x5E, 0x0D, 0x2B, 0x07, 0x5A, 0x12, 0x75, 0x5B,
	0x58, 0x02, 0x09, 0x0C, 0x02, 0x4A, 0x5A, 0x04, 0x2C, 0x2B, 0x13, 0x19,
	0x0E, 0x0A, 0x05, 0x4A, 0x41, 0x0F, 0x2D, 0x18, 0x15, 0x07, 0x13, 0x36,
	0x0A, 0x13, 0x5B, 0x05, 0x71, 0x0A, 0x19, 0x06, 0x0A, 0x3B, 0x03, 0x52,
	0x5B, 0x3A, 0x26, 0x3C, 0x1B, 0x1A, 0x3C, 0x2D, 0x08, 0x03, 0x1F, 0x33,
	0x2C, 0x5B, 0x50, 0x04, 0x0F, 0x31, 0x1D, 0x31, 0x1A, 0x33, 0x33, 0x38,
	0x54, 0x56, 0x39, 0x1B, 0x2A, 0x16, 0x57, 0x3F, 0x06, 0x59, 0x0B, 0x23,
	0x59, 0x69, 0x01, 0x36, 0x23, 0x2D, 0x31, 0x15, 0x3B, 0x3A, 0x22, 0x2C,
	0x0F, 0x51, 0x2D, 0x29, 0x2B, 0x47, 0x17, 0x0B, 0x12, 0x14, 0x21, 0x25,
	0x06, 0x44, 0x18, 0x3B, 0x2D, 0x00, 0x18, 0x70, 0x09, 0x34, 0x22, 0x18,
	0x2E, 0x5F, 0x57, 0x23, 0x5E, 0x75, 0x5E, 0x0C, 0x5D, 0x2D, 0x71, 0x05,
	0x55, 0x0A, 0x13, 0x74, 0x22, 0x36, 0x16, 0x20, 0x25, 0x5A, 0x05, 0x37,
	0x5D, 0x16, 0x01, 0x0D, 0x0C, 0x2E, 0x32, 0x2D, 0x4A, 0x34, 0x28, 0x11,
	0x04, 0x4E, 0x5B, 0x23, 0x32, 0x5B, 0x25, 0x0D, 0x1D, 0x37, 0x43, 0x37,
	0x14, 0x23, 0x25, 0x5B, 0x2B, 0x38, 0x5E, 0x2E, 0x54, 0x14, 0x01, 0x19,
	0x18, 0x09, 0x38, 0x28, 0x05, 0x70, 0x0F, 0x00, 0x2C, 0x44, 0x2A, 0x19,
	0x0B, 0x07, 0x58, 0x76, 0x2A, 0x0F, 0x05, 0x5A, 0x13, 0x5A, 0x19, 0x39,
	0x3C, 0x27, 0x2D, 0x53, 0x45, 0x26, 0x38, 0x59, 0x56, 0x3C, 0x1B, 0x2C,
	0x2F, 0x53, 0x01, 0x44, 0x01, 0x1D, 0x10, 0x07, 0x1F, 0x20, 0x54, 0x36,
	0x1A, 0x27, 0x70, 0x1E, 0x35, 0x20, 0x00, 0x10, 0x36, 0x0D, 0x1D, 0x5F,
	0x20, 0x29, 0x0C, 0x18, 0x5B, 0x3A, 0x02, 0x1B, 0x05, 0x1C, 0x2D, 0x5D,
	0x31, 0x3E, 0x1D, 0x36, 0x39, 0x02, 0x02, 0x0F, 0x15, 0x1F, 0x08, 0x0F,
	0x32, 0x3A, 0x3A, 0x39, 0x1A, 0x44, 0x00, 0x27, 0x55, 0x34, 0x5F, 0x34,
	0x15, 0x58, 0x16, 0x44, 0x7B, 0x1D, 0x24, 0x3B, 0x19, 0x10, 0x3E, 0x09,
	0x1D, 0x5F, 0x1B, 0x43, 0x05, 0x3D, 0x59, 0x2B, 0x20, 0x2C, 0x2D, 0x59,
	0x28, 0x0E, 0x10, 0x08, 0x3D, 0x24, 0x3E, 0x55, 0x00, 0x3B, 0x24, 0x25,
	0x51, 0x29, 0x58, 0x30, 0x05, 0x4A, 0x59, 0x1C, 0x74, 0x43, 0x12, 0x56,
	0x02, 0x20, 0x14, 0x37, 0x38, 0x2F, 0x2E, 0x34, 0x4A, 0x39, 0x05, 0x34,
	0x1B, 0x05, 0x1E, 0x3F, 0x28, 0x55, 0x57, 0x0B, 0x11, 0x2A, 0x5F, 0x15,
	0x5A, 0x3F, 0x34, 0x3A, 0x10, 0x00, 0x27, 0x03, 0x14, 0x36, 0x0A, 0x5A,
	0x0D, 0x3A, 0x2C, 0x0A, 0x03, 0x16, 0x19, 0x26, 0x03, 0x5B, 0x71, 0x36,
	0x2C, 0x36, 0x3D, 0x36, 0x34, 0x36, 0x18, 0x31, 0x2A, 0x54, 0x14, 0x3E,
	0x1B, 0x34, 0x59, 0x3B, 0x2D, 0x58, 0x35, 0x5B, 0x38, 0x04, 0x06, 0x3B,
	0x36, 0x52, 0x06, 0x00, 0x3A, 0x2E, 0x35, 0x2A, 0x33, 0x1B, 0x2B, 0x31,
	0x24, 0x1B, 0x27, 0x23, 0x4A, 0x22, 0x23, 0x73, 0x34, 0x34, 0x20, 0x1C,
	0x1B, 0x18, 0x06, 0x27, 0x0A, 0x75, 0x54, 0x4A, 0x1C, 0x32, 0x7B, 0x08,
	0x04, 0x01, 0x5A, 0x76, 0x00, 0x4E, 0x34, 0x00, 0x73, 0x1F, 0x26, 0x5C,
	0x1B, 0x73, 0x5B, 0x0D, 0x41, 0x13, 0x3A, 0x0F, 0x4A, 0x45, 0x33, 0x7A,
	0x24, 0x08, 0x41, 0x06, 0x75, 0x19, 0x31, 0x22, 0x58, 0x7B, 0x47, 0x00,
	0x59, 0x24, 0x17, 0x14, 0x19, 0x45, 0x5E, 0x3A, 0x3E, 0x35, 0x59, 0x2F,
	0x23, 0x5D, 0x29, 0x04, 0x3A, 0x09, 0x01, 0x0C, 0x04, 0x31, 0x75, 0x34,
	0x12, 0x3C, 0x24, 0x71, 0x0E, 0x0B, 0x56, 0x18, 0x37, 0x23, 0x14, 0x5B,
	0x20, 0x06, 0x02, 0x4E, 0x5E, 0x0F, 0x11, 0x0A, 0x26, 0x14, 0x58, 0x73,
	0x34, 0x0D, 0x1E, 0x3B, 0x15, 0x5B, 0x3B, 0x05, 0x00, 0x37, 0x0A, 0x51,
	0x00, 0x20, 0x01, 0x5C, 0x26, 0x01, 0x1D, 0x2A, 0x02, 0x08, 0x1B, 0x2C,
	0x30, 0x26, 0x14, 0x16, 0x04, 0x2E, 0x38, 0x27, 0x1D, 0x5B, 0x24, 0x5C,
	0x08, 0x57, 0x3C, 0x75, 0x27, 0x30, 0x5D, 0x2F, 0x28, 0x58, 0x14, 0x0C,
	0x07, 0x37, 0x14, 0x13, 0x39, 0x2F, 0x2E, 0x54, 0x18, 0x37, 0x59, 0x03,
	0x0B, 0x24, 0x56, 0x5D, 0x33, 0x0F, 0x2F, 0x5D, 0x40, 0x06, 0x3A, 0x02,
	0x29, 0x53, 0x7B, 0x5F, 0x26, 0x22, 0x5D, 0x28, 0x58, 0x37, 0x2A, 0x04,
	0x2A, 0x36, 0x2A, 0x08, 0x1C, 0x35, 0x0E, 0x55, 0x14, 0x1F, 0x26, 0x0D,
	0x15, 0x59, 0x21, 0x70, 0x3B, 0x2E, 0x09, 0x20, 0x0A, 0x35, 0x51, 0x2A,
	0x3F, 0x69, 0x35, 0x31, 0x0B, 0x11, 0x74, 0x04, 0x11, 0x17, 0x5C, 0x26,
	0x0A, 0x02, 0x25, 0x1C, 0x72, 0x0A, 0x17, 0x5E, 0x1D, 0x24, 0x08, 0x03,
	0x39, 0x1C, 0x75, 0x0E, 0x39, 0x22, 0x2D, 0x2E, 0x3B, 0x34, 0x5D, 0x26,
	0x00, 0x58, 0x4E, 0x0C, 0x03, 0x1A, 0x0F, 0x4A, 0x5F, 0x09, 0x7A, 0x43,
	0x57, 0x39, 0x2D, 0x76, 0x0D, 0x05, 0x0A, 0x31, 0x75, 0x59, 0x11, 0x34,
	0x23, 0x30, 0x1E, 0x25, 0x5D, 0x5C, 0x31, 0x1F, 0x17, 0x16, 0x27, 0x2A,
	0x35, 0x3B, 0x27, 0x3A, 0x26, 0x1A, 0x2D, 0x14, 0x23, 0x28, 0x23, 0x31,
	0x19, 0x3B, 0x70, 0x0E, 0x53, 0x07, 0x0E, 0x0F, 0x0E, 0x39, 0x28, 0x0D,
	0x15, 0x55, 0x31, 0x0F, 0x3B, 0x2D, 0x1C, 0x54, 0x19, 0x27, 0x72, 0x58,
	0x35, 0x0D, 0x13, 0x32, 0x08, 0x22, 0x57, 0x59, 0x26, 0x55, 0x18, 0x56,
	0x5E, 0x27, 0x0D, 0x20, 0x14, 0x5B, 0x0A, 0x19, 0x02, 0x39, 0x31, 0x0A,
	0x0F, 0x50, 0x18, 0x24, 0x05, 0x1E, 0x0E, 0x26, 0x18, 0x20, 0x5B, 0x31,
	0x00, 0x5C, 0x2F, 0x1D, 0x53, 0x37, 0x5B, 0x70, 0x19, 0x04, 0x5D, 0x1C,
	0x3A, 0x07, 0x39, 0x0C, 0x58, 0x12, 0x0B, 0x53, 0x5F, 0x0C, 0x36, 0x27,
	0x4E, 0x3B, 0x3D, 0x37, 0x0F, 0x18, 0x39, 0x11, 0x24, 0x3A, 0x05, 0x3C,
	0x0D, 0x0C, 0x15, 0x04, 0x5B, 0x06, 0x73, 0x0E, 0x58, 0x0A, 0x5A, 0x0C,
	0x5C, 0x57, 0x5D, 0x2E, 0x0D, 0x01, 0x10, 0x18, 0x09, 0x27, 0x5D, 0x2F,
	0x5F, 0x5E, 0x17, 0x14, 0x14, 0x37, 0x26, 0x05, 0x36, 0x10, 0x5B, 0x11,
	0x30, 0x0E, 0x37, 0x5A, 0x19, 0x69, 0x02, 0x3B, 0x00, 0x24, 0x0A, 0x1D,
	0x03, 0x03, 0x1A, 0x77, 0x58, 0x32, 0x08, 0x27, 0x3A, 0x36, 0x34, 0x57,
	0x20, 0x2B, 0x20, 0x34, 0x41, 0x03, 0x20, 0x19, 0x0C, 0x1D, 0x04, 0x2D,
	0x21, 0x54, 0x5A, 0x1E, 0x37, 0x09, 0x19, 0x17, 0x31, 0x09, 0x20, 0x13,
	0x3A, 0x19, 0x3A, 0x14, 0x12, 0x3F, 0x18, 0x75, 0x0D, 0x10, 0x04, 0x5E,
	0x04, 0x0A, 0x58, 0x2B, 0x07, 0x3B, 0x1A, 0x29, 0x2A, 0x27, 0x09, 0x09,
	0x04, 0x28, 0x02, 0x75, 0x22, 0x2F, 0x00, 0x06, 0x38, 0x2D, 0x54, 0x20,
	0x44, 0x0D, 0x26, 0x12, 0x56, 0x24, 0x07, 0x1F, 0x37, 0x45, 0x1F, 0x25,
	0x06, 0x03, 0x20, 0x31, 0x73, 0x35, 0x53, 0x3C, 0x00, 0x73, 0x47, 0x39,
	0x21, 0x5C, 0x0F, 0x3B, 0x57, 0x3E, 0x20, 0x69, 0x1A, 0x55, 0x1A, 0x13,
	0x38, 0x1D, 0x03, 0x0A, 0x2C, 0x24, 0x22, 0x0B, 0x5E, 0x2A, 0x06, 0x02,
	0x55, 0x26, 0x5A, 0x15, 0x2A, 0x30, 0x03, 0x09, 0x1A, 0x06, 0x17, 0x57,
	0x3D, 0x10, 0x2B, 0x11, 0x5C, 0x0A, 0x37, 0x1F, 0x18, 0x1F, 0x06, 0x29,
	0x27, 0x38, 0x0B, 0x58, 0x23, 0x5D, 0x36, 0x24, 0x3E, 0x7A, 0x3C, 0x11,
	0x03, 0x23, 0x73, 0x5B, 0x24, 0x05, 0x24, 0x26, 0x0A, 0x2B, 0x0C, 0x1D,
	0x33, 0x28, 0x0B, 0x0A, 0x59, 0x7A, 0x38, 0x11, 0x17, 0x1A, 0x12, 0x03,
	0x0B, 0x37, 0x5F, 0x7B, 0x02, 0x0B, 0x01, 0x59, 0x34, 0x08, 0x0B, 0x45,
	0x18, 0x29, 0x36, 0x17, 0x04, 0x40, 0x12, 0x2D, 0x35, 0x3A, 0x1E, 0x70,
	0x27, 0x33, 0x41, 0x20, 0x26, 0x1B, 0x19, 0x18, 0x01, 0x1B, 0x59, 0x00,
	0x20, 0x08, 0x6D, 0x0A, 0x02, 0x3B, 0x1D, 0x6D, 0x04, 0x4E, 0x0D, 0x27,
	0x2A, 0x0E, 0x10, 0x21, 0x59, 0x36, 0x0A, 0x12, 0x28, 0x44, 0x69, 0x25,
	0x14, 0x21, 0x3B, 0x25, 0x19, 0x07, 0x03, 0x01, 0x6D, 0x5C, 0x4E, 0x0F,
	0x39, 0x2D, 0x0F, 0x0D, 0x5A, 0x0E, 0x0F, 0x02, 0x2D, 0x1C, 0x06, 0x26,
	0x5B, 0x07, 0x2F, 0x40, 0x20, 0x26, 0x29, 0x1B, 0x1A, 0x17, 0x54, 0x04,
	0x2A, 0x1E, 0x12, 0x19, 0x52, 0x20, 0x44, 0x07, 0x01, 0x34, 0x0A, 0x5A,
	0x27, 0x3C, 0x2A, 0x01, 0x1B, 0x77, 0x01, 0x11, 0x14, 0x11, 0x14, 0x5B,
	0x3B, 0x0D, 0x1A, 0x0A, 0x59, 0x2A, 0x3F, 0x3D, 0x09, 0x47, 0x19, 0x36,
	0x24, 0x21, 0x43, 0x15, 0x5C, 0x59, 0x09, 0x39, 0x38, 0x04, 0x52, 0x3B,
	0x24, 0x17, 0x56, 0x1B, 0x24, 0x0E, 0x14, 0x57, 0x44, 0x20, 0x0E, 0x04,
	0x1E, 0x3D, 0x29, 0x58, 0x55, 0x5A, 0x0F, 0x26, 0x3A, 0x23, 0x2A, 0x07,
	0x77, 0x3C, 0x2B, 0x38, 0x5E, 0x69, 0x5D, 0x18, 0x38, 0x0F, 0x12, 0x0E,
	0x05, 0x41, 0x3C, 0x21, 0x0E, 0x1B, 0x0B, 0x2C, 0x30, 0x5B, 0x2F, 0x05,
	0x5C, 0x6D, 0x1F, 0x55, 0x21, 0x5F, 0x0C, 0x3C, 0x0A, 0x41, 0x3A, 0x30,
	0x20, 0x20, 0x08, 0x31, 0x71, 0x0D, 0x14, 0x1D, 0x5A, 0x2F, 0x01, 0x00,
	0x56, 0x0F, 0x74, 0x5E, 0x58, 0x05, 0x33, 0x23, 0x5C, 0x1B, 0x02, 0x44,
	0x2C, 0x0E, 0x25, 0x20, 0x3B, 0x07, 0x20, 0x17, 0x0B, 0x40, 0x34, 0x3D,
	0x35, 0x20, 0x18, 0x00, 0x5B, 0x2E, 0x2D, 0x0E, 0x0D, 0x55, 0x13, 0x2D,
	0x09, 0x26, 0x5F, 0x32, 0x04, 0x25, 0x75, 0x1A, 0x26, 0x29, 0x1F, 0x33,
	0x01, 0x19, 0x2A, 0x03, 0x12, 0x5E, 0x55, 0x5C, 0x3E, 0x70, 0x1E, 0x35,
	0x0F, 0x5D, 0x36, 0x20, 0x16, 0x0C, 0x28, 0x31, 0x43, 0x35, 0x0F, 0x3D,
	0x0D, 0x19, 0x4A, 0x45, 0x2F, 0x28, 0x2B, 0x00, 0x0F, 0x19, 0x0C, 0x26,
	0x59, 0x5C, 0x3B, 0x36, 0x54, 0x07, 0x1A, 0x26, 0x05, 0x5B, 0x31, 0x29,
	0x24, 0x08, 0x39, 0x0D, 0x3A, 0x1C, 0x73, 0x1F, 0x56, 0x20, 0x52, 0x69,
	0x0D, 0x1B, 0x3D, 0x44, 0x7A, 0x08, 0x22, 0x58, 0x0D, 0x09, 0x28, 0x15,
	0x19, 0x5E, 0x09, 0x0F, 0x13, 0x0A, 0x0A, 0x23, 0x58, 0x00, 0x0B, 0x0E,
	0x1A, 0x36, 0x51, 0x09, 0x1F, 0x0D, 0x0E, 0x11, 0x22, 0x28, 0x37, 0x55,
	0x31, 0x0D, 0x19, 0x20, 0x47, 0x15, 0x03, 0x3F, 0x28, 0x5E, 0x12, 0x41,
	0x5D, 0x15, 0x18, 0x38, 0x26, 0x40, 0x75, 0x16, 0x3B, 0x08, 0x40, 0x1A,
	0x19, 0x1B, 0x0B, 0x2C, 0x38, 0x18, 0x58, 0x14, 0x27, 0x37, 0x5B, 0x13,
	0x59, 0x19, 0x14, 0x28, 0x39, 0x16, 0x09, 0x38, 0x2A, 0x0D, 0x1C, 0x1E,
	0x2C, 0x16, 0x06, 0x5E, 0x0A, 0x34, 0x01, 0x11, 0x26, 0x23, 0x33, 0x0F,
	0x59, 0x57, 0x29, 0x36, 0x19, 0x53, 0x3F, 0x3F, 0x2B, 0x02, 0x17, 0x09,
	0x3A, 0x6D, 0x34, 0x53, 0x21, 0x07, 0x3A, 0x15, 0x0B, 0x22, 0x00, 0x72,
	0x3E, 0x31, 0x1A, 0x01, 0x3A, 0x0A, 0x10, 0x5A, 0x03, 0x76, 0x19, 0x26,
	0x0B, 0x21, 0x73, 0x1C, 0x22, 0x07, 0x06, 0x21, 0x15, 0x09, 0x5B, 0x02,
	0x10, 0x5A, 0x50, 0x5A, 0x0A, 0x2B, 0x21, 0x03, 0x23, 0x1A, 0x10, 0x54,
	0x0E, 0x02, 0x0D, 0x24, 0x39, 0x54, 0x14, 0x3B, 0x25, 0x16, 0x53, 0x04,
	0x07, 0x2D, 0x5A, 0x34, 0x18, 0x0A, 0x35, 0x09, 0x17, 0x21, 0x01, 0x1B,
	0x2E, 0x50, 0x5C, 0x23, 0x75, 0x34, 0x2C, 0x29, 0x5E, 0x6D, 0x5A, 0x0E,
	0x56, 0x39, 0x75, 0x5F, 0x2B, 0x00, 0x19, 0x35, 0x5D, 0x16, 0x1A, 0x1B,
	0x24, 0x14, 0x17, 0x28, 0x52, 0x2A, 0x54, 0x59, 0x22, 0x00, 0x26, 0x03,
	0x27, 0x2A, 0x58, 0x37, 0x24, 0x57, 0x1D, 0x0E, 0x77, 0x16, 0x56, 0x08,
	0x52, 0x3B, 0x54, 0x55, 0x0C, 0x26, 0x14, 0x1B, 0x0F, 0x0C, 0x40, 0x71,
	0x43, 0x12, 0x24, 0x5B, 0x09, 0x47, 0x57, 0x37, 0x18, 0x0C, 0x2D, 0x25,
	0x1A, 0x29, 0x01, 0x1E, 0x58, 0x41, 0x06, 0x01, 0x29, 0x3B, 0x38, 0x0A,
	0x3A, 0x00, 0x00, 0x08, 0x0A, 0x2F, 0x1F, 0x02, 0x18, 0x2F, 0x70, 0x0A,
	0x36, 0x2C, 0x5C, 0x14, 0x3B, 0x0F, 0x5E, 0x5F, 0x32, 0x3B, 0x57, 0x36,
	0x5E, 0x23, 0x20, 0x12, 0x01, 0x1A, 0x0A, 0x04, 0x00, 0x41, 0x26, 0x31,
	0x24, 0x16, 0x14, 0x00, 0x34, 0x2E, 0x39, 0x1B, 0x52, 0x75, 0x23, 0x51,
	0x56, 0x5A, 0x08, 0x5B, 0x2C, 0x0C, 0x24, 0x0F, 0x36, 0x0B, 0x02, 0x1C,
	0x33, 0x0F, 0x10, 0x1C, 0x25, 0x23, 0x5A, 0x52, 0x2C, 0x5E, 0x17, 0x2A,
	0x34, 0x20, 0x52, 0x0D, 0x24, 0x07, 0x1C, 0x33, 0x0B, 0x2A, 0x07, 0x1F,
	0x1F, 0x16, 0x02, 0x2D, 0x2C, 0x06, 0x13, 0x3C, 0x12, 0x1C, 0x03, 0x77,
	0x25, 0x29, 0x2C, 0x1E, 0x25, 0x43, 0x14, 0x09, 0x1C, 0x6D, 0x0A, 0x31,
	0x1C, 0x24, 0x04, 0x1A, 0x34, 0x3C, 0x5F, 0x72, 0x18, 0x22, 0x04, 0x0F,
	0x32, 0x2B, 0x3B, 0x29, 0x44, 0x21, 0x2E, 0x20, 0x21, 0x52, 0x32, 0x0F,
	0x0D, 0x5E, 0x05, 0x0E, 0x2E, 0x53, 0x34, 0x40, 0x23, 0x2B, 0x10, 0x0F,
	0x26, 0x0B, 0x0B, 0x1B, 0x3B, 0x2F, 0x3A, 0x5F, 0x3B, 0x41, 0x24, 0x2D,
	0x3A, 0x52, 0x37, 0x2F, 0x23, 0x0D, 0x1B, 0x0A, 0x12, 0x71, 0x0F, 0x38,
	0x08, 0x27, 0x24, 0x0B, 0x2F, 0x5F, 0x04, 0x7A, 0x06, 0x15, 0x5B, 0x5D,
	0x38, 0x1D, 0x2D, 0x03, 0x1C, 0x27, 0x2A, 0x11, 0x04, 0x26, 0x2A, 0x59,
	0x27, 0x1F, 0x1E, 0x15, 0x16, 0x2D, 0x03, 0x1A, 0x26, 0x02, 0x32, 0x0D,
	0x13, 0x18, 0x5A, 0x29, 0x04, 0x0D, 0x35, 0x1F, 0x0C, 0x5A, 0x2E, 0x15,
	0x24, 0x4E, 0x08, 0x07, 0x24, 0x38, 0x11, 0x16, 0x53, 0x32, 0x5F, 0x54,
	0x1F, 0x53, 0x0C, 0x06, 0x4A, 0x17, 0x08, 0x2E, 0x24, 0x1B, 0x0A, 0x44,
	0x05, 0x5E, 0x58, 0x5E, 0x53, 0x0D, 0x2F, 0x09, 0x29, 0x0E, 0x18, 0x06,
	0x0F, 0x57, 0x40, 0x34, 0x3C, 0x25, 0x1D, 0x00, 0x71, 0x3C, 0x1B, 0x23,
	0x03, 0x2A, 0x47, 0x58, 0x0C, 0x1E, 0x28, 0x5F, 0x2F, 0x38, 0x44, 0x18,
	0x59, 0x18, 0x22, 0x3F, 0x38, 0x43, 0x07, 0x28, 0x0C, 0x01, 0x0F, 0x58,
	0x5F, 0x2D, 0x16, 0x38, 0x37, 0x45, 0x1C, 0x20, 0x07, 0x31, 0x28, 0x24,
	0x33, 0x5C, 0x0D, 0x5A, 0x19, 0x2C, 0x28, 0x20, 0x09, 0x24, 0x30, 0x1F,
	0x06, 0x23, 0x23, 0x1A, 0x2D, 0x06, 0x0B, 0x2E, 0x32, 0x1C, 0x3B, 0x00,
	0x23, 0x0C, 0x21, 0x53, 0x29, 0x2D, 0x06, 0x39, 0x2F, 0x2B, 0x3E, 0x6D,
	0x1A, 0x14, 0x2C, 0x29, 0x24, 0x58, 0x04, 0x0A, 0x3B, 0x71, 0x15, 0x0C,
	0x24, 0x06, 0x71, 0x1C, 0x03, 0x5C, 0x07, 0x69, 0x5C, 0x04, 0x00, 0x12,
	0x26, 0x29, 0x27, 0x41, 0x19, 0x11, 0x15, 0x4E, 0x08, 0x01, 0x36, 0x08,
	0x33, 0x41, 0x3F, 0x12, 0x02, 0x0F, 0x5E, 0x5A, 0x0D, 0x23, 0x00, 0x1C,
	0x3C, 0x34, 0x54, 0x31, 0x58, 0x5B, 0x18, 0x58, 0x56, 0x08, 0x03, 0x70,
	0x1A, 0x05, 0x45, 0x39, 0x2E, 0x3D, 0x55, 0x41, 0x53, 0x75, 0x47, 0x12,
	0x58, 0x0D, 0x27, 0x18, 0x33, 0x56, 0x58, 0x12, 0x5E, 0x17, 0x00, 0x1B,
	0x6D, 0x0E, 0x54, 0x18, 0x13, 0x3B, 0x55, 0x0D, 0x07, 0x1B, 0x38, 0x5A,
	0x39, 0x3A, 0x02, 0x27, 0x19, 0x17, 0x59, 0x1F, 0x27, 0x27, 0x18, 0x08,
	0x0A, 0x0D, 0x2B, 0x28, 0x07, 0x38, 0x7B, 0x1F, 0x2D, 0x57, 0x22, 0x0A,
	0x5F, 0x52, 0x0B, 0x32, 0x18, 0x0A, 0x3B, 0x06, 0x22, 0x24, 0x5F, 0x2F,
	0x26, 0x18, 0x37, 0x5D, 0x34, 0x5C, 0x18, 0x11, 0x5A, 0x2A, 0x20, 0x28,
	0x2A, 0x25, 0x57, 0x36, 0x5D, 0x35, 0x0A, 0x35, 0x5F, 0x58, 0x36, 0x3A,
	0x1B, 0x03, 0x5B, 0x17, 0x0A, 0x25, 0x27, 0x5C, 0x27, 0x23, 0x0A, 0x5C,
	0x3B, 0x7A, 0x47, 0x10, 0x5C, 0x02, 0x3A, 0x1D, 0x19, 0x57, 0x11, 0x11,
	0x0F, 0x11, 0x26, 0x2E, 0x75, 0x20, 0x54, 0x37, 0x0A, 0x69, 0x26, 0x07,
	0x36, 0x5D, 0x0E, 0x21, 0x33, 0x00, 0x2C, 0x38, 0x34, 0x56, 0x08, 0x26,
	0x75, 0x5E, 0x04, 0x03, 0x25, 0x75, 0x26, 0x39, 0x3A, 0x11, 0x6D, 0x38,
	0x37, 0x58, 0x31, 0x01, 0x5B, 0x09, 0x3A, 0x52, 0x2E, 0x39, 0x36, 0x26,
	0x3F, 0x0F, 0x09, 0x31, 0x45, 0x0E, 0x0A, 0x16, 0x11, 0x26, 0x59, 0x23,
	0x27, 0x03, 0x1D, 0x53, 0x35, 0x35, 0x37, 0x58, 0x02, 0x15, 0x34, 0x57,
	0x19, 0x01, 0x0D, 0x58, 0x13, 0x38, 0x5D, 0x36, 0x1C, 0x4A, 0x03, 0x39,
	0x77, 0x2A, 0x15, 0x08, 0x29, 0x14, 0x01, 0x31, 0x45, 0x52, 0x18, 0x58,
	0x17, 0x25, 0x52, 0x77, 0x22, 0x36, 0x38, 0x05, 0x1A, 0x47, 0x07, 0x2B,
	0x08, 0x17, 0x03, 0x19, 0x07, 0x58, 0x12, 0x5B, 0x07, 0x04, 0x05, 0x35,
	0x2B, 0x2F, 0x41, 0x13, 0x35, 0x20, 0x07, 0x18, 0x40, 0x77, 0x01, 0x14,
	0x22, 0x0C, 0x20, 0x5E, 0x2E, 0x00, 0x58, 0x0A, 0x1D, 0x3B, 0x17, 0x0D,
	0x77, 0x16, 0x14, 0x01, 0x1A, 0x21, 0x43, 0x14, 0x5F, 0x0F, 0x21, 0x5E,
	0x13, 0x19, 0x01, 0x24, 0x5C, 0x2C, 0x08, 0x32, 0x34, 0x1F, 0x4A, 0x03,
	0x40, 0x11, 0x47, 0x54, 0x08, 0x38, 0x23, 0x3C, 0x07, 0x38, 0x20, 0x74,
	0x59, 0x3B, 0x06, 0x09, 0x2C, 0x5B, 0x11, 0x0A, 0x5B, 0x73, 0x08, 0x27,
	0x36, 0x20, 0x06, 0x5C, 0x53, 0x0A, 0x3F, 0x38, 0x3B, 0x0D, 0x5D, 0x31,
	0x2E, 0x1D, 0x14, 0x57, 0x1A, 0x3A, 0x59, 0x57, 0x0B, 0x5D, 0x3B, 0x23,
	0x36, 0x20, 0x32, 0x75, 0x1B, 0x32, 0x3A, 0x5A, 0x69, 0x5D, 0x31, 0x08,
	0x5E, 0x0C, 0x5B, 0x56, 0x24, 0x5F, 0x24, 0x43, 0x2A, 0x26, 0x2C, 0x70,
	0x5A, 0x50, 0x5E, 0x5A, 0x69, 0x3C, 0x20, 0x2D, 0x52, 0x38, 0x08, 0x07,
	0x0B, 0x58, 0x73, 0x5B, 0x52, 0x0B, 0x09, 0x0E, 0x3C, 0x0F, 0x39, 0x59,
	0x14, 0x55, 0x53, 0x37, 0x09, 0x3B, 0x18, 0x57, 0x22, 0x0A, 0x34, 0x1F,
	0x11, 0x38, 0x5A, 0x10, 0x47, 0x03, 0x39, 0x12, 0x1B, 0x01, 0x18, 0x18,
	0x1D, 0x3B, 0x36, 0x54, 0x1D, 0x40, 0x7B, 0x58, 0x36, 0x08, 0x3A, 0x33,
	0x47, 0x03, 0x07, 0x18, 0x2E, 0x59, 0x29, 0x1D, 0x19, 0x17, 0x07, 0x25,
	0x41, 0x08, 0x38, 0x58, 0x38, 0x41, 0x09, 0x0A, 0x38, 0x29, 0x3C, 0x0E,
	0x32, 0x23, 0x50, 0x20, 0x19, 0x01, 0x58, 0x1B, 0x56, 0x3F, 0x09, 0x0E,
	0x2E, 0x39, 0x03, 0x74, 0x5A, 0x0C, 0x07, 0x3F, 0x77, 0x27, 0x37, 0x0B,
	0x22, 0x69, 0x1D, 0x03, 0x0B, 0x1B, 0x31, 0x0F, 0x22, 0x1B, 0x2F, 0x0B,
	0x18, 0x20, 0x25, 0x0D, 0x05, 0x54, 0x05, 0x3A, 0x39, 0x73, 0x43, 0x2E,
	0x0C, 0x1F, 0x2A, 0x1E, 0x52, 0x23, 0x5F, 0x0C, 0x5E, 0x07, 0x03, 0x02,
	0x32, 0x21, 0x23, 0x5A, 0x1A, 0x21, 0x34, 0x26, 0x5C, 0x0A, 0x69, 0x19,
	0x23, 0x06, 0x03, 0x12, 0x20, 0x0F, 0x5D, 0x21, 0x24, 0x38, 0x15, 0x2D,
	0x58, 0x6D, 0x06, 0x1B, 0x0A, 0x0F, 0x73, 0x3E, 0x17, 0x3C, 0x11, 0x34,
	0x55, 0x19, 0x14, 0x02, 0x26, 0x5C, 0x07, 0x20, 0x20, 0x05, 0x59, 0x1B,
	0x14, 0x40, 0x2B, 0x1E, 0x0B, 0x58, 0x5C, 0x30, 0x5B, 0x14, 0x26, 0x58,
	0x28, 0x24, 0x57, 0x03, 0x2D, 0x06, 0x24, 0x15, 0x1B, 0x3C, 0x24, 0x3C,
	0x23, 0x5D, 0x59, 0x34, 0x0E, 0x0D, 0x00, 0x0E, 0x33, 0x18, 0x10, 0x14,
	0x0A, 0x0D, 0x55, 0x26, 0x45, 0x1E, 0x12, 0x47, 0x50, 0x5D, 0x18, 0x31,
	0x23, 0x03, 0x06, 0x40, 0x37, 0x0F, 0x17, 0x1F, 0x5A, 0x16, 0x5D, 0x53,
	0x08, 0x2A, 0x29, 0x14, 0x0C, 0x02, 0x40, 0x17, 0x5D, 0x0C, 0x3E, 0x2A,
	0x69, 0x0D, 0x03, 0x59, 0x1C, 0x33, 0x3B, 0x2E, 0x3E, 0x3F, 0x0B, 0x5F,
	0x25, 0x28, 0x04, 0x21, 0x23, 0x37, 0x34, 0x06, 0x7B, 0x3C, 0x00, 0x09,
	0x3C, 0x18, 0x5A, 0x14, 0x5E, 0x3A, 0x15, 0x06, 0x25, 0x5F, 0x44, 0x70,
	0x0A, 0x03, 0x5C, 0x1F, 0x37, 0x55, 0x20, 0x01, 0x5C, 0x30, 0x15, 0x0D,
	0x14, 0x39, 0x16, 0x18, 0x23, 0x2D, 0x25, 0x30, 0x28, 0x3B, 0x5D, 0x28,
	0x0B, 0x0E, 0x14, 0x1A, 0x01, 0x07, 0x5A, 0x12, 0x03, 0x58, 0x11, 0x14,
	0x4E, 0x5B, 0x12, 0x12, 0x04, 0x0A, 0x1D, 0x3B, 0x06, 0x20, 0x13, 0x34,
	0x24, 0x6D, 0x19, 0x51, 0x5A, 0x08, 0x00, 0x25, 0x13, 0x0F, 0x02, 0x34,
	0x1E, 0x2F, 0x03, 0x2C, 0x14, 0x3A, 0x12, 0x0C, 0x0F, 0x26, 0x07, 0x00,
	0x3B, 0x32, 0x20, 0x3B, 0x13, 0x16, 0x53, 0x0B, 0x09, 0x15, 0x5C, 0x00,
	0x05, 0x1B, 0x03, 0x1B, 0x38, 0x16, 0x59, 0x32, 0x45, 0x0D, 0x33, 0x00,
	0x30, 0x0B, 0x0A, 0x0A, 0x3D, 0x58, 0x56, 0x59, 0x11, 0x3D, 0x55, 0x0F,
	0x2F, 0x0E, 0x2F, 0x2A, 0x36, 0x5A, 0x13, 0x5E, 0x07, 0x24, 0x1A, 0x00,
	0x47, 0x54, 0x0C, 0x59, 0x73, 0x5E, 0x0E, 0x22, 0x39, 0x3A, 0x07, 0x12,
	0x00, 0x27, 0x0A, 0x39, 0x30, 0x02, 0x3C, 0x71, 0x04, 0x59, 0x26, 0x52,
	0x73, 0x3D, 0x00, 0x03, 0x06, 0x18, 0x1F, 0x04, 0x58, 0x0F, 0x37, 0x5C,
	0x37, 0x5F, 0x58, 0x0B, 0x55, 0x58, 0x17, 0x03, 0x12, 0x47, 0x3B, 0x3D,
	0x1C, 0x30, 0x1D, 0x27, 0x3D, 0x58, 0x0E, 0x5C, 0x25, 0x0A, 0x39, 0x24,
	0x2E, 0x2F, 0x41, 0x33, 0x7B, 0x55, 0x34, 0x18, 0x5B, 0x70, 0x02, 0x00,
	0x41, 0x0D, 0x70, 0x00, 0x0D, 0x18, 0x5F, 0x73, 0x20, 0x55, 0x23, 0x3B,
	0x2B, 0x0A, 0x50, 0x18, 0x5D, 0x26, 0x5E, 0x54, 0x24, 0x20, 0x33, 0x3E,
	0x35, 0x02, 0x1E, 0x34, 0x22, 0x1B, 0x06, 0x2A, 0x34, 0x2B, 0x13, 0x14,
	0x12, 0x2B, 0x15, 0x58, 0x5F, 0x53, 0x30, 0x1E, 0x04, 0x1D, 0x5C, 0x1B,
	0x58, 0x57, 0x01, 0x05, 0x15, 0x3E, 0x36, 0x0D, 0x1D, 0x6D, 0x1D, 0x25,
	0x05, 0x03, 0x75, 0x28, 0x15, 0x1D, 0x29, 0x3B, 0x3F, 0x07, 0x09, 0x3D,
	0x71, 0x35, 0x19, 0x3A, 0x2D, 0x70, 0x0E, 0x0E, 0x45, 0x12, 0x75, 0x3A,
	0x27, 0x0D, 0x18, 0x7A, 0x2B, 0x0F, 0x3A, 0x38, 0x29, 0x02, 0x35, 0x18,
	0x27, 0x32, 0x5D, 0x39, 0x56, 0x07, 0x16, 0x20, 0x37, 0x18, 0x0E, 0x3A,
	0x0B, 0x38, 0x5B, 0x27, 0x71, 0x5D, 0x15, 0x1A, 0x1F, 0x0B, 0x3C, 0x52,
	0x41, 0x1B, 0x2D, 0x5F, 0x59, 0x1B, 0x2E, 0x18, 0x3B, 0x0B, 0x41, 0x59,
	0x37, 0x19, 0x0F, 0x0C, 0x27, 0x31, 0x5E, 0x0D, 0x26, 0x3A, 0x25, 0x47,
	0x12, 0x21, 0x22, 0x1B, 0x20, 0x54, 0x34, 0x3C, 0x69, 0x08, 0x07, 0x00,
	0x13, 0x76, 0x01, 0x19, 0x5B, 0x19, 0x13, 0x5B, 0x09, 0x5A, 0x0A, 0x07,
	0x38, 0x06, 0x57, 0x53, 0x33, 0x43, 0x2F, 0x5B, 0x52, 0x31, 0x23, 0x58,
	0x28, 0x20, 0x70, 0x06, 0x2E, 0x03, 0x58, 0x06, 0x38, 0x2C, 0x0F, 0x07,
	0x0C, 0x59, 0x03, 0x1F, 0x0D, 0x0E, 0x21, 0x50, 0x22, 0x21, 0x2B, 0x59,
	0x31, 0x3B, 0x1C, 0x2C, 0x5B, 0x17, 0x03, 0x39, 0x30, 0x59, 0x0E, 0x59,
	0x0E, 0x37, 0x02, 0x12, 0x23, 0x0D, 0x71, 0x47, 0x0B, 0x3C, 0x0D, 0x7B,
	0x38, 0x31, 0x18, 0x5B, 0x09, 0x2A, 0x17, 0x0C, 0x2F, 0x71, 0x1C, 0x56,
	0x1A, 0x0D, 0x6D, 0x3B, 0x52, 0x5F, 0x0D, 0x17, 0x2B, 0x0B, 0x1E, 0x2D,
	0x15, 0x58, 0x2F, 0x03, 0x5D, 0x11, 0x2F, 0x4A, 0x14, 0x0F, 0x00, 0x3B,
	0x51, 0x58, 0x21, 0x20, 0x5F, 0x11, 0x07, 0x18, 0x32, 0x5A, 0x52, 0x0A,
	0x0D, 0x12, 0x02, 0x53, 0x05, 0x38, 0x7B, 0x5F, 0x15, 0x0C, 0x11, 0x70,
	0x36, 0x1B, 0x45, 0x1A, 0x28, 0x08, 0x4A, 0x05, 0x0F, 0x27, 0x02, 0x35,
	0x19, 0x2C, 0x2C, 0x19, 0x1B, 0x17, 0x0F, 0x32, 0x3C, 0x04, 0x17, 0x1D,
	0x74, 0x38, 0x19, 0x5D, 0x1C, 0x71, 0x2D, 0x15, 0x5F, 0x1D, 0x16, 0x5D,
	0x55, 0x5E, 0x0E, 0x72, 0x1D, 0x26, 0x06, 0x1F, 0x37, 0x2E, 0x2A, 0x17,
	0x5A, 0x3B, 0x2B, 0x18, 0x3F, 0x0D, 0x0C, 0x0D, 0x55, 0x0A, 0x24, 0x13,
	0x5C, 0x0E, 0x06, 0x3D, 0x2F, 0x00, 0x14, 0x3D, 0x1C, 0x6D, 0x05, 0x34,
	0x00, 0x2D, 0x16, 0x22, 0x37, 0x5A, 0x08, 0x70, 0x3A, 0x37, 0x19, 0x52,
	0x74, 0x5A, 0x23, 0x1E, 0x20, 0x0E, 0x00, 0x37, 0x1B, 0x2E, 0x69, 0x5D,
	0x39, 0x0D, 0x24, 0x12, 0x18, 0x18, 0x3E, 0x31, 0x17, 0x1D, 0x37, 0x21,
	0x32, 0x69, 0x3A, 0x56, 0x0D, 0x39, 0x28, 0x08, 0x03, 0x37, 0x23, 0x05,
	0x0B, 0x11, 0x0B, 0x5B, 0x03, 0x58, 0x57, 0x00, 0x21, 0x70, 0x06, 0x0E,
	0x57, 0x03, 0x26, 0x54, 0x13, 0x02, 0x07, 0x2F, 0x1D, 0x39, 0x26, 0x5C,
	0x35, 0x27, 0x05, 0x5B, 0x11, 0x30, 0x1F, 0x4A, 0x1F, 0x23, 0x7A, 0x5A,
	0x53, 0x1C, 0x40, 0x29, 0x0A, 0x4A, 0x2B, 0x1B, 0x7B, 0x34, 0x0C, 0x22,
	0x1B, 0x05, 0x00, 0x32, 0x21, 0x5C, 0x05, 0x5A, 0x51, 0x3E, 0x40, 0x24,
	0x2F, 0x31, 0x1F, 0x0C, 0x11, 0x3C, 0x37, 0x25, 0x12, 0x28, 0x18, 0x00,
	0x1D, 0x29, 0x2E, 0x08, 0x07, 0x3A, 0x52, 0x14, 0x23, 0x0F, 0x36, 0x33,
	0x32, 0x3E, 0x00, 0x5F, 0x1E, 0x05, 0x19, 0x17, 0x34, 0x24, 0x6D, 0x3B,
	0x29, 0x5F, 0x2F, 0x20, 0x0F, 0x53, 0x0B, 0x2A, 0x76, 0x5B, 0x0B, 0x1E,
	0x13, 0x15, 0x1E, 0x56, 0x2C, 0x5D, 0x37, 0x39, 0x25, 0x34, 0x00, 0x76,
	0x39, 0x08, 0x5E, 0x1E, 0x09, 0x01, 0x31, 0x07, 0x53, 0x1A, 0x59, 0x26,
	0x0F, 0x02, 0x12, 0x55, 0x0B, 0x59, 0x40, 0x69, 0x54, 0x2A, 0x24, 0x31,
	0x26, 0x09, 0x17, 0x5F, 0x53, 0x3B, 0x22, 0x1B, 0x1A, 0x27, 0x23, 0x1E,
	0x1B, 0x1C, 0x12, 0x1A, 0x0F, 0x39, 0x3E, 0x0E, 0x00, 0x1C, 0x29, 0x1F,
	0x59, 0x2B, 0x08, 0x17, 0x59, 0x06, 0x7A, 0x23, 0x58, 0x38, 0x2C, 0x14,
	0x19, 0x35, 0x5C, 0x58, 0x71, 0x0E, 0x33, 0x3E, 0x3E, 0x73, 0x3B, 0x53,
	0x19, 0x3B, 0x10, 0x28, 0x10, 0x39, 0x3C, 0x28, 0x2F, 0x10, 0x0F, 0x5C,
	0x75, 0x14, 0x31, 0x02, 0x5D, 0x06, 0x03, 0x37, 0x5C, 0x0F, 0x10, 0x28,
	0x4E, 0x0F, 0x44, 0x0A, 0x36, 0x00, 0x1C, 0x22, 0x18, 0x3C, 0x2E, 0x05,
	0x3C, 0x6D, 0x0D, 0x55, 0x1F, 0x2F, 0x25, 0x5A, 0x52, 0x1E, 0x58, 0x3A,
	0x16, 0x51, 0x2F, 0x07, 0x2E, 0x08, 0x2D, 0x39, 0x0E, 0x1A, 0x54, 0x3B,
	0x0F, 0x0D, 0x77, 0x22, 0x0F, 0x36, 0x03, 0x21, 0x2B, 0x2A, 0x37, 0x58,
	0x24, 0x2D, 0x0D, 0x5F, 0x3D, 0x36, 0x26, 0x55, 0x0C, 0x40, 0x0A, 0x05,
	0x33, 0x21, 0x1B, 0x36, 0x18, 0x59, 0x3D, 0x44, 0x18, 0x59, 0x18, 0x19,
	0x1B, 0x29, 0x5A, 0x19, 0x02, 0x05, 0x2D, 0x5E, 0x39, 0x3E, 0x12, 0x2B,
	0x0A, 0x26, 0x26, 0x59, 0x06, 0x3C, 0x12, 0x1A, 0x0A, 0x2F, 0x09, 0x34,
	0x59, 0x59, 0x75, 0x16, 0x25, 0x3E, 0x3E, 0x15, 0x3A, 0x08, 0x04, 0x1D,
	0x2C, 0x1C, 0x34, 0x56, 0x2A, 0x2A, 0x1F, 0x4E, 0x3C, 0x01, 0x29, 0x5E,
	0x2A, 0x45, 0x11, 0x3B, 0x1F, 0x12, 0x27, 0x29, 0x3B, 0x04, 0x39, 0x23,
	0x33, 0x32, 0x3C, 0x0B, 0x0C, 0x25, 0x7B, 0x3D, 0x4A, 0x29, 0x1F, 0x71,
	0x1F, 0x07, 0x0B, 0x53, 0x30, 0x5A, 0x2B, 0x3B, 0x3B, 0x38, 0x43, 0x54,
	0x27, 0x1D, 0x18, 0x38, 0x22, 0x39, 0x33, 0x2E, 0x1E, 0x32, 0x3B, 0x01,
	0x12, 0x1E, 0x59, 0x21, 0x1B, 0x27, 0x14, 0x54, 0x45, 0x25, 0x01, 0x04,
	0x35, 0x39, 0x21, 0x01, 0x47, 0x03, 0x2D, 0x3B, 0x14, 0x0A, 0x2E, 0x38,
	0x52, 0x73, 0x38, 0x2B, 0x0F, 0x06, 0x75, 0x5E, 0x08, 0x01, 0x3C, 0x3A,
	0x09, 0x54, 0x3C, 0x5B, 0x2C, 0x04, 0x36, 0x08, 0x40, 0x7A, 0x08, 0x18,
	0x1D, 0x1F, 0x0E, 0x2B, 0x17, 0x1F, 0x05, 0x09, 0x07, 0x0F, 0x41, 0x53,
	0x2E, 0x0A, 0x0E, 0x39, 0x03, 0x26, 0x09, 0x13, 0x00, 0x0F, 0x10, 0x3A,
	0x12, 0x1C, 0x3E, 0x75, 0x1A, 0x29, 0x41, 0x11, 0x2A, 0x38, 0x15, 0x5A,
	0x5C, 0x0B, 0x09, 0x53, 0x29, 0x01, 0x12, 0x19, 0x33, 0x18, 0x11, 0x10,
	0x1C, 0x16, 0x36, 0x24, 0x38, 0x54, 0x51, 0x00, 0x5F, 0x17, 0x5B, 0x33,
	0x23, 0x44, 0x32, 0x5B, 0x02, 0x01, 0x0D, 0x2A, 0x36, 0x4E, 0x3D, 0x04,
	0x72, 0x15, 0x4A, 0x45, 0x04, 0x69, 0x20, 0x11, 0x3E, 0x1A, 0x76, 0x1E,
	0x09, 0x02, 0x3D, 0x21, 0x1B, 0x51, 0x3A, 0x24, 0x04, 0x19, 0x07, 0x21,
	0x52, 0x14, 0x05, 0x2B, 0x14, 0x0D, 0x31, 0x3F, 0x54, 0x1C, 0x04, 0x74,
	0x20, 0x16, 0x36, 0x3F, 0x12, 0x19, 0x59, 0x57, 0x5A, 0x12, 0x05, 0x03,
	0x3E, 0x0F, 0x1B, 0x0B, 0x2F, 0x0D, 0x07, 0x30, 0x18, 0x27, 0x3E, 0x2D,
	0x26, 0x1A, 0x58, 0x23, 0x5F, 0x3A, 0x18, 0x37, 0x37, 0x0F, 0x2B, 0x3D,
	0x54, 0x57, 0x06, 0x11, 0x22, 0x29, 0x5E, 0x26, 0x37, 0x43, 0x03, 0x2B,
	0x58, 0x03, 0x0F, 0x00, 0x03, 0x1D, 0x35, 0x09, 0x50, 0x24, 0x0F, 0x37,
	0x2F, 0x1B, 0x3F, 0x5F, 0x3A, 0x54, 0x0B, 0x5E, 0x3A, 0x6D, 0x28, 0x03,
	0x24, 0x27, 0x1A, 0x43, 0x39, 0x56, 0x01, 0x09, 0x54, 0x58, 0x41, 0x1B,
	0x37, 0x1F, 0x06, 0x37, 0x23, 0x24, 0x19, 0x36, 0x2B, 0x5A, 0x33, 0x58,
	0x08, 0x5D, 0x07, 0x31, 0x05, 0x0B, 0x3D, 0x52, 0x7B, 0x38, 0x53, 0x27,
	0x2D, 0x16, 0x5B, 0x05, 0x3B, 0x2E, 0x0E, 0x16, 0x0A, 0x58, 0x04, 0x11,
	0x54, 0x22, 0x25, 0x1B, 0x01, 0x3E, 0x10, 0x3D, 0x3E, 0x09, 0x01, 0x13,
	0x09, 0x1A, 0x28, 0x0E, 0x56, 0x0C, 0x2E, 0x08, 0x2D, 0x03, 0x14, 0x25,
	0x01, 0x28, 0x08, 0x22, 0x33, 0x06, 0x5A, 0x02, 0x0F, 0x22, 0x35, 0x3E,
	0x22, 0x5D, 0x13, 0x07, 0x35, 0x07, 0x36, 0x5D, 0x10, 0x24, 0x1B, 0x1E,
	0x19, 0x18, 0x58, 0x38, 0x1D, 0x08, 0x06, 0x34, 0x27, 0x17, 0x26, 0x15,
	0x47, 0x31, 0x3F, 0x13, 0x1B, 0x03, 0x24, 0x3E, 0x13, 0x23, 0x55, 0x07,
	0x5C, 0x2A, 0x34, 0x2B, 0x16, 0x19, 0x3E, 0x69, 0x2B, 0x20, 0x56, 0x33,
	0x69, 0x24, 0x11, 0x09, 0x13, 0x03, 0x26, 0x07, 0x26, 0x5F, 0x3A, 0x35,
	0x55, 0x20, 0x3B, 0x06, 0x05, 0x20, 0x3B, 0x40, 0x07, 0x25, 0x59, 0x39,
	0x40, 0x0A, 0x1C, 0x0B, 0x16, 0x2A, 0x09, 0x0A, 0x29, 0x05, 0x32, 0x37,
	0x54, 0x26, 0x26, 0x2E, 0x03, 0x00, 0x58, 0x18, 0x01, 0x04, 0x06, 0x06,
	0x5E, 0x12, 0x72, 0x01, 0x27, 0x18, 0x02, 0x0F, 0x5A, 0x2C, 0x3F, 0x28,
	0x1A, 0x5A, 0x4A, 0x28, 0x07, 0x15, 0x05, 0x23, 0x3A, 0x44, 0x27, 0x25,
	0x24, 0x5F, 0x19, 0x25, 0x21, 0x52, 0x17, 0x29, 0x2D, 0x1B, 0x34, 0x45,
	0x2E, 0x38, 0x18, 0x08, 0x09, 0x3E, 0x69, 0x5F, 0x06, 0x28, 0x01, 0x25,
	0x21, 0x56, 0x14, 0x09, 0x25, 0x04, 0x03, 0x5A, 0x3F, 0x0F, 0x27, 0x2B,
	0x2C, 0x3F, 0x74, 0x16, 0x4E, 0x3A, 0x58, 0x13, 0x2D, 0x11, 0x57, 0x29,
	0x03, 0x1E, 0x29, 0x2F, 0x31, 0x77, 0x14, 0x29, 0x22, 0x3B, 0x01, 0x36,
	0x25, 0x07, 0x2E, 0x15, 0x47, 0x20, 0x19, 0x24, 0x12, 0x39, 0x38, 0x22,
	0x0D, 0x0F, 0x0E, 0x2B, 0x16, 0x2A, 0x09, 0x0A, 0x10, 0x3D, 0x06, 0x3A,
	0x1B, 0x2A, 0x0B, 0x0D, 0x13, 0x05, 0x1B, 0x19, 0x52, 0x16, 0x16, 0x50,
	0x28, 0x5A, 0x30, 0x0B, 0x57, 0x41, 0x1D, 0x2E, 0x23, 0x37, 0x1C, 0x0C,
	0x72, 0x16, 0x4A, 0x37, 0x0C, 0x00, 0x0E, 0x55, 0x0B, 0x01, 0x38, 0x26,
	0x30, 0x19, 0x1F, 0x7A, 0x0A, 0x02, 0x1E, 0x23, 0x07, 0x3D, 0x15, 0x56,
	0x00, 0x76, 0x0B, 0x27, 0x18, 0x03, 0x75, 0x0D, 0x19, 0x2F, 0x21, 0x24,
	0x24, 0x1B, 0x00, 0x03, 0x2F, 0x43, 0x4E, 0x2A, 0x0F, 0x76, 0x24, 0x14,
	0x0F, 0x44, 0x30, 0x18, 0x52, 0x0D, 0x27, 0x26, 0x5E, 0x17, 0x28, 0x0D,
	0x74, 0x3F, 0x14, 0x57, 0x1E, 0x37, 0x0E, 0x07, 0x5D, 0x28, 0x70, 0x54,
	0x33, 0x5F, 0x5B, 0x04, 0x04, 0x00, 0x1A, 0x22, 0x74, 0x23, 0x50, 0x20,
	0x3B, 0x0F, 0x54, 0x08, 0x37, 0x3D, 0x2A, 0x29, 0x2B, 0x2C, 0x09, 0x2F,
	0x24, 0x57, 0x02, 0x22, 0x1A, 0x59, 0x19, 0x29, 0x13, 0x08, 0x09, 0x32,
	0x1D, 0x2F, 0x2B, 0x0E, 0x36, 0x2A, 0x06, 0x37, 0x26, 0x2C, 0x20, 0x19,
	0x11, 0x0A, 0x06, 0x36, 0x28, 0x20, 0x5D, 0x29, 0x2B, 0x3B, 0x03, 0x5C,
	0x22, 0x0A, 0x0E, 0x11, 0x47, 0x05, 0x5A, 0x0C, 0x2D, 0x0D, 0x0A, 0x3E,
	0x2A, 0x10, 0x5D, 0x28, 0x39, 0x24, 0x3B, 0x1A, 0x58, 0x23, 0x0D, 0x34,
	0x2A, 0x07, 0x57, 0x44, 0x69, 0x5E, 0x36, 0x03, 0x21, 0x74, 0x35, 0x0C,
	0x24, 0x08, 0x17, 0x20, 0x55, 0x1E, 0x25, 0x38, 0x24, 0x00, 0x14, 0x1F,
	0x20, 0x36, 0x28, 0x14, 0x26, 0x75, 0x24, 0x55, 0x0B, 0x2F, 0x76, 0x02,
	0x2F, 0x38, 0x5B, 0x25, 0x59, 0x31, 0x2A, 0x01, 0x17, 0x43, 0x0B, 0x1D,
	0x27, 0x07, 0x59, 0x59, 0x21, 0x01, 0x27, 0x2A, 0x23, 0x5C, 0x20, 0x16,
	0x23, 0x03, 0x45, 0x20, 0x75, 0x43, 0x56, 0x04, 0x28, 0x16, 0x16, 0x0E,
	0x25, 0x0E, 0x2F, 0x36, 0x29, 0x2A, 0x1A, 0x1A, 0x26, 0x57, 0x3A, 0x11,
	0x31, 0x06, 0x0D, 0x0D, 0x3F, 0x28, 0x27, 0x2A, 0x2B, 0x5D, 0x10, 0x3C,
	0x54, 0x1A, 0x29, 0x77, 0x27, 0x39, 0x3C, 0x03, 0x24, 0x06, 0x00, 0x26,
	0x05, 0x2B, 0x5A, 0x06, 0x5C, 0x13, 0x07, 0x1C, 0x53, 0x3D, 0x29, 0x32,
	0x21, 0x0D, 0x5D, 0x22, 0x03, 0x47, 0x58, 0x19, 0x00, 0x69, 0x01, 0x02,
	0x3E, 0x2E, 0x74, 0x3F, 0x32, 0x23, 0x03, 0x0D, 0x16, 0x2E, 0x3C, 0x0C,
	0x29, 0x38, 0x16, 0x0B, 0x3B, 0x1B, 0x1A, 0x2F, 0x14, 0x0A, 0x24, 0x16,
	0x04, 0x3D, 0x2A, 0x28, 0x2D, 0x34, 0x0D, 0x04, 0x35, 0x2E, 0x09, 0x5B,
	0x38, 0x18, 0x07, 0x08, 0x3F, 0x3F, 0x33, 0x3C, 0x32, 0x45, 0x0E, 0x38,
	0x19, 0x00, 0x05, 0x08, 0x03, 0x36, 0x53, 0x36, 0x1C, 0x69, 0x2A, 0x0F,
	0x1D, 0x19, 0x0F, 0x5B, 0x51, 0x00, 0x27, 0x29, 0x27, 0x30, 0x3C, 0x32,
	0x2D, 0x2A, 0x59, 0x56, 0x20, 0x38, 0x3D, 0x16, 0x3E, 0x02, 0x01, 0x25,
	0x19, 0x37, 0x2F, 0x69, 0x1D, 0x20, 0x06, 0x2C, 0x24, 0x2F, 0x20, 0x04,
	0x26, 0x2B, 0x35, 0x59, 0x25, 0x21, 0x0B, 0x3E, 0x55, 0x16, 0x3B, 0x32,
	0x14, 0x59, 0x3F, 0x12, 0x0D, 0x24, 0x16, 0x1B, 0x21, 0x7B, 0x3C, 0x33,
	0x2F, 0x0F, 0x17, 0x59, 0x0A, 0x2D, 0x24, 0x0F, 0x58, 0x00, 0x0D, 0x27,
	0x0D, 0x38, 0x27, 0x1D, 0x32, 0x14, 0x25, 0x00, 0x28, 0x18, 0x03, 0x3B,
	0x12, 0x04, 0x3B, 0x32, 0x24, 0x25, 0x58, 0x0D, 0x3A, 0x5A, 0x04, 0x00,
	0x08, 0x69, 0x01, 0x23, 0x08, 0x1B, 0x25, 0x2B, 0x0A, 0x38, 0x52, 0x2D,
	0x3B, 0x29, 0x16, 0x04, 0x11, 0x20, 0x18, 0x3E, 0x09, 0x70, 0x04, 0x55,
	0x24, 0x2F, 0x23, 0x21, 0x0F, 0x1D, 0x39, 0x0E, 0x59, 0x0F, 0x04, 0x3A,
	0x31, 0x3F, 0x23, 0x1B, 0x2F, 0x28, 0x1F, 0x1B, 0x26, 0x3D, 0x13, 0x05,
	0x31, 0x37, 0x1F, 0x06, 0x38, 0x4A, 0x26, 0x13, 0x31, 0x55, 0x09, 0x2D,
	0x40, 0x11, 0x22, 0x07, 0x0A, 0x01, 0x0B, 0x55, 0x2E, 0x1E, 0x5B, 0x34,
	0x2A, 0x2D, 0x2B, 0x11, 0x24, 0x38, 0x28, 0x14, 0x0E, 0x17, 0x00, 0x51,
	0x3E, 0x00, 0x21, 0x0B, 0x18, 0x06, 0x39, 0x70, 0x25, 0x2B, 0x14, 0x2C,
	0x1B, 0x3B, 0x04, 0x2A, 0x12, 0x2B, 0x39, 0x2B, 0x2B, 0x08, 0x75, 0x0B,
	0x27, 0x45, 0x03, 0x0A, 0x06, 0x53, 0x26, 0x11, 0x37, 0x09, 0x0F, 0x0D,
	0x3D, 0x03, 0x55, 0x57, 0x1F, 0x2E, 0x25, 0x25, 0x2A, 0x34, 0x09, 0x04,
	0x15, 0x04, 0x22, 0x13, 0x7A, 0x47, 0x0F, 0x39, 0x0F, 0x01, 0x29, 0x4E,
	0x26, 0x53, 0x10, 0x28, 0x38, 0x1C, 0x2D, 0x2A, 0x36, 0x0C, 0x19, 0x03,
	0x00, 0x47, 0x30, 0x5D, 0x38, 0x21, 0x3D, 0x23, 0x3A, 0x31, 0x08, 0x21,
	0x3B, 0x5C, 0x0D, 0x3A, 0x3E, 0x27, 0x19, 0x03, 0x71, 0x08, 0x28, 0x07,
	0x26, 0x77, 0x01, 0x04, 0x03, 0x28, 0x6D, 0x07, 0x22, 0x25, 0x13, 0x31,
	0x0E, 0x26, 0x19, 0x3A, 0x70, 0x1F, 0x06, 0x45, 0x31, 0x25, 0x03, 0x58,
	0x25, 0x31, 0x0D, 0x34, 0x0C, 0x2F, 0x02, 0x23, 0x21, 0x2B, 0x05, 0x1E,
	0x07, 0x20, 0x2A, 0x3A, 0x26, 0x30, 0x2E, 0x02, 0x39, 0x2D, 0x69, 0x35,
	0x0C, 0x3B, 0x28, 0x1B, 0x16, 0x20, 0x23, 0x07, 0x07, 0x39, 0x53, 0x2C,
	0x3C, 0x1B, 0x05, 0x26, 0x01, 0x19, 0x7B, 0x47, 0x0F, 0x09, 0x03, 0x2D,
	0x27, 0x22, 0x24, 0x3A, 0x0B, 0x25, 0x0C, 0x36, 0x07, 0x21, 0x5C, 0x35,
	0x09, 0x29, 0x21, 0x14, 0x24, 0x3A, 0x0E, 0x08, 0x00, 0x54, 0x05, 0x21,
	0x0F, 0x29, 0x04, 0x1A, 0x13, 0x10, 0x0E, 0x18, 0x1D, 0x1F, 0x09, 0x38,
	0x38, 0x3E, 0x26, 0x2C, 0x38, 0x06, 0x3C, 0x13, 0x26, 0x29, 0x20, 0x2D,
	0x02, 0x70, 0x15, 0x28, 0x3E, 0x2F, 0x31, 0x5B, 0x0C, 0x5C, 0x52, 0x06,
	0x18, 0x59, 0x09, 0x3E, 0x07, 0x39, 0x06, 0x2C, 0x44, 0x03, 0x3E, 0x36,
	0x29, 0x03, 0x73, 0x00, 0x06, 0x45, 0x1B, 0x2F, 0x54, 0x0D, 0x22, 0x07,
	0x18, 0x35, 0x2F, 0x08, 0x39, 0x72, 0x1C, 0x20, 0x0B, 0x2E, 0x11, 0x08,
	0x19, 0x2B, 0x12, 0x03, 0x0E, 0x36, 0x37, 0x5D, 0x33, 0x01, 0x30, 0x25,
	0x0A, 0x2A, 0x28, 0x20, 0x09, 0x0E, 0x2C, 0x2D, 0x0A, 0x56, 0x5A, 0x06,
	0x34, 0x06, 0x26, 0x5D, 0x2A, 0x23, 0x0F, 0x3E, 0x22, 0x15, 0x07, 0x22,
	0x25, 0x3A, 0x16, 0x35, 0x06, 0x2D, 0x26, 0x13, 0x1C, 0x2E, 0x0A, 0x1C,
	0x0F, 0x1A, 0x31, 0x1E, 0x06, 0x15, 0x14, 0x4A, 0x25, 0x0C, 0x26, 0x07,
	0x16, 0x05, 0x1D, 0x09, 0x1F, 0x2A, 0x26, 0x3F, 0x0B, 0x09, 0x26, 0x24,
	0x2C, 0x06, 0x36, 0x39, 0x3A, 0x00, 0x14, 0x2D, 0x4A, 0x06, 0x2C, 0x1B,
	0x1A, 0x18, 0x09, 0x5C, 0x0F, 0x14, 0x53, 0x3C, 0x1F, 0x0C, 0x21, 0x2D,
	0x57, 0x2C, 0x10, 0x23, 0x33, 0x16, 0x1B, 0x1B, 0x2B, 0x55, 0x1A, 0x18,
	0x69, 0x0A, 0x07, 0x3D, 0x44, 0x77, 0x15, 0x04, 0x3D, 0x24, 0x27, 0x38,
	0x18, 0x21, 0x32, 0x2F, 0x54, 0x53, 0x2C, 0x5C, 0x03, 0x06, 0x13, 0x14,
	0x18, 0x30, 0x22, 0x23, 0x24, 0x09, 0x0E, 0x35, 0x4E, 0x2F, 0x1C, 0x1B,
	0x36, 0x10, 0x0D, 0x2A, 0x75, 0x2E, 0x27, 0x1E, 0x18, 0x25, 0x3D, 0x28,
	0x0D, 0x2A, 0x04, 0x59, 0x53, 0x2B, 0x22, 0x2A, 0x26, 0x18, 0x1D, 0x09,
	0x17, 0x2F, 0x4E, 0x34, 0x28, 0x2A, 0x39, 0x37, 0x16, 0x29, 0x15, 0x25,
	0x34, 0x02, 0x27, 0x11, 0x07, 0x58, 0x27, 0x5E, 0x2D, 0x24, 0x27, 0x24,
	0x3F, 0x2D, 0x2E, 0x34, 0x58, 0x26, 0x76, 0x58, 0x06, 0x36, 0x13, 0x0D,
	0x0E, 0x15, 0x0A, 0x22, 0x0D, 0x1C, 0x17, 0x3E, 0x31, 0x69, 0x08, 0x25,
	0x27, 0x18, 0x0D, 0x54, 0x2E, 0x34, 0x06, 0x21, 0x20, 0x2B, 0x2D, 0x2D,
	0x13, 0x25, 0x54, 0x41, 0x31, 0x38, 0x58, 0x2D, 0x3B, 0x23, 0x10, 0x2F,
	0x35, 0x02, 0x5F, 0x70, 0x3D, 0x2B, 0x0B, 0x00, 0x27, 0x16, 0x54, 0x0A,
	0x1C, 0x17, 0x19, 0x20, 0x04, 0x44, 0x25, 0x54, 0x2C, 0x00, 0x53, 0x3B,
	0x1B, 0x50, 0x26, 0x1B, 0x34, 0x1C, 0x50, 0x1F, 0x3A, 0x06, 0x3F, 0x3B,
	0x00, 0x28, 0x70, 0x38, 0x2F, 0x3A, 0x2F, 0x6D, 0x08, 0x20, 0x28, 0x00,
	0x04, 0x2A, 0x23, 0x20, 0x3A, 0x06, 0x35, 0x4A, 0x24, 0x12, 0x2F, 0x38,
	0x0F, 0x34, 0x5E, 0x04, 0x04, 0x57, 0x5E, 0x04, 0x03, 0x2E, 0x0F, 0x19,
	0x26, 0x30, 0x1C, 0x36, 0x29, 0x12, 0x03, 0x3A, 0x25, 0x27, 0x03, 0x01,
	0x21, 0x22, 0x0C, 0x1A, 0x73, 0x3F, 0x0C, 0x34, 0x1D, 0x04, 0x16, 0x30,
	0x19, 0x3E, 0x10, 0x54, 0x31, 0x1F, 0x1C, 0x71, 0x00, 0x23, 0x5E, 0x0E,
	0x10, 0x28, 0x36, 0x5A, 0x3A, 0x2C, 0x58, 0x57, 0x16, 0x28, 0x27, 0x0F,
	0x0A, 0x5B, 0x38, 0x24, 0x2E, 0x2A, 0x3F, 0x26, 0x2B, 0x20, 0x32, 0x28,
	0x2F, 0x35, 0x3E, 0x2B, 0x08, 0x25, 0x2A, 0x5D, 0x13, 0x3C, 0x3E, 0x2D,
	0x15, 0x27, 0x2B, 0x38, 0x07, 0x03, 0x53, 0x29, 0x5D, 0x08, 0x3C, 0x37,
	0x3B, 0x3A, 0x2A, 0x36, 0x22, 0x17, 0x3F, 0x0B, 0x35, 0x31, 0x03, 0x44,
	0x32, 0x07, 0x02, 0x1F, 0x19, 0x0A, 0x34, 0x52, 0x1A, 0x5E, 0x0B, 0x3A,
	0x03, 0x5A, 0x3C, 0x03, 0x16, 0x11, 0x3E, 0x25, 0x16, 0x07, 0x2A, 0x57,
	0x1D, 0x2E, 0x21, 0x18, 0x3D, 0x2C, 0x0F, 0x3E, 0x50, 0x5B, 0x19, 0x31,
	0x47, 0x26, 0x28, 0x53, 0x2C, 0x04, 0x23, 0x5C, 0x28, 0x1B, 0x20, 0x29,
	0x3E, 0x0A, 0x00, 0x35, 0x06, 0x0A, 0x27, 0x00, 0x07, 0x53, 0x58, 0x33,
	0x18, 0x16, 0x27, 0x29, 0x5F, 0x75, 0x0F, 0x2B, 0x2F, 0x3A, 0x1A, 0x59,
	0x16, 0x00, 0x13, 0x74, 0x35, 0x0B, 0x1F, 0x0C, 0x05, 0x26, 0x04, 0x3F,
	0x0C, 0x0A, 0x3E, 0x33, 0x20, 0x1A, 0x0B, 0x38, 0x56, 0x2F, 0x03, 0x7A,
	0x34, 0x09, 0x0F, 0x1A, 0x13, 0x28, 0x2B, 0x25, 0x07, 0x21, 0x5D, 0x2E,
	0x3C, 0x32, 0x71, 0x07, 0x27, 0x19, 0x40, 0x3A, 0x05, 0x23, 0x08, 0x1C,
	0x31, 0x0B, 0x22, 0x57, 0x2E, 0x36, 0x01, 0x0E, 0x1F, 0x5F, 0x0D, 0x47,
	0x22, 0x00, 0x5C, 0x05, 0x20, 0x52, 0x59, 0x20, 0x0E, 0x25, 0x25, 0x22,
	0x2A, 0x23, 0x58, 0x2E, 0x1B, 0x26, 0x6D, 0x3C, 0x22, 0x0A, 0x0E, 0x2E,
	0x5F, 0x14, 0x02, 0x08, 0x0B, 0x21, 0x06, 0x03, 0x2E, 0x7B, 0x14, 0x2E,
	0x05, 0x2F, 0x27, 0x08, 0x0C, 0x56, 0x3B, 0x0E, 0x16, 0x28, 0x26, 0x25,
	0x11, 0x20, 0x2A, 0x45, 0x27, 0x3B, 0x3E, 0x25, 0x29, 0x02, 0x21, 0x55,
	0x2F, 0x3B, 0x59, 0x0B, 0x5C, 0x26, 0x22, 0x05, 0x03, 0x2B, 0x18, 0x06,
	0x28, 0x12, 0x2F, 0x06, 0x06, 0x58, 0x0F, 0x3F, 0x33, 0x0B, 0x06, 0x03,
	0x23, 0x10, 0x3C, 0x08, 0x03, 0x2F, 0x35, 0x24, 0x3F, 0x10, 0x09, 0x0C,
	0x5E, 0x0A, 0x71, 0x55, 0x06, 0x5D, 0x5A, 0x05, 0x21, 0x04, 0x24, 0x52,
	0x24, 0x0A, 0x19, 0x29, 0x13, 0x13, 0x09, 0x26, 0x45, 0x5F, 0x13, 0x14,
	0x08, 0x36, 0x13, 0x13, 0x5A, 0x16, 0x2A, 0x2C, 0x25, 0x27, 0x51, 0x20,
	0x3C, 0x76, 0x1F, 0x25, 0x0F, 0x26, 0x2B, 0x04, 0x22, 0x5D, 0x22, 0x77,
	0x02, 0x26, 0x19, 0x0C, 0x74, 0x00, 0x2B, 0x1D, 0x26, 0x2F, 0x5D, 0x20,
	0x3C, 0x07, 0x01, 0x05, 0x04, 0x3B, 0x20, 0x11, 0x27, 0x56, 0x37, 0x1B,
	0x00, 0x24, 0x26, 0x1A, 0x39, 0x13, 0x25, 0x2E, 0x5A, 0x00, 0x16, 0x2D,
	0x24, 0x0D, 0x00, 0x15, 0x2A, 0x0D, 0x2A, 0x02, 0x07, 0x08, 0x16, 0x01,
	0x07, 0x35, 0x0A, 0x51, 0x27, 0x3A, 0x2D, 0x2B, 0x54, 0x3F, 0x05, 0x16,
	0x23, 0x29, 0x14, 0x3E, 0x29, 0x35, 0x2A, 0x17, 0x18, 0x28, 0x06, 0x2B,
	0x58, 0x32, 0x03, 0x35, 0x30, 0x2D, 0x38, 0x13, 0x5B, 0x20, 0x06, 0x20,
	0x14, 0x38, 0x25, 0x5A, 0x3E, 0x08, 0x3E, 0x0B, 0x2C, 0x5E, 0x69, 0x3E,
	0x39, 0x2B, 0x44, 0x0B, 0x03, 0x54, 0x3A, 0x24, 0x26, 0x2F, 0x24, 0x5B,
	0x08, 0x04, 0x0B, 0x29, 0x5B, 0x5D, 0x1A, 0x14, 0x4A, 0x2B, 0x27, 0x20,
	0x38, 0x23, 0x58, 0x0C, 0x17, 0x34, 0x2A, 0x58, 0x2A, 0x0F, 0x0B, 0x56,
	0x2A, 0x1B, 0x31, 0x3C, 0x22, 0x34, 0x0A, 0x18, 0x16, 0x12, 0x5C, 0x2A,
	0x1A, 0x3D, 0x2A, 0x27, 0x22, 0x1B, 0x5D, 0x4E, 0x5B, 0x59, 0x12, 0x22,
	0x54, 0x59, 0x28, 0x16, 0x54, 0x4A, 0x03, 0x2E, 0x37, 0x29, 0x32, 0x5B,
	0x21, 0x26, 0x18, 0x22, 0x0C, 0x2F, 0x30, 0x00, 0x33, 0x03, 0x3A, 0x03,
	0x3B, 0x0E, 0x26, 0x25, 0x77, 0x15, 0x06, 0x27, 0x3A, 0x0E, 0x35, 0x33,
	0x02, 0x2D, 0x6D, 0x26, 0x0E, 0x26, 0x33, 0x11, 0x04, 0x03, 0x2C, 0x24,
	0x08, 0x22, 0x0F, 0x45, 0x58, 0x20, 0x2A, 0x28, 0x3B, 0x05, 0x16, 0x1D,
	0x00, 0x28, 0x2D, 0x21, 0x5C, 0x2C, 0x0A, 0x29, 0x29, 0x0D, 0x30, 0x0D,
	0x5D, 0x36, 0x0E, 0x0D, 0x23, 0x25, 0x01, 0x1A, 0x23, 0x25, 0x22, 0x31,
	0x38, 0x0C, 0x3F, 0x0A, 0x10, 0x29, 0x59, 0x45, 0x24, 0x25, 0x22, 0x2B,
	0x22, 0x29, 0x03, 0x26, 0x16, 0x28, 0x28, 0x27, 0x28, 0x28, 0x3F, 0x5A,
	0x0E, 0x14, 0x14, 0x22, 0x22, 0x03, 0x26, 0x0A, 0x27, 0x03, 0x25, 0x00,
	0x54, 0x57, 0x07, 0x24, 0x1A, 0x28, 0x5D, 0x2D, 0x21, 0x22, 0x2D, 0x5B,
	0x02, 0x2E, 0x2A, 0x16, 0x1A, 0x22, 0x28, 0x28, 0x1B, 0x5B, 0x0E, 0x12,
	0x0B, 0x10, 0x09, 0x40, 0x2D, 0x25, 0x53, 0x3A, 0x5D, 0x14, 0x16, 0x30,
	0x21, 0x3A, 0x1A, 0x59, 0x30, 0x23, 0x39, 0x2C, 0x2D, 0x00, 0x14, 0x3A,
	0x13, 0x23, 0x0C, 0x04, 0x00, 0x09, 0x23, 0x4A, 0x0C, 0x25, 0x06, 0x09,
	0x59, 0x03, 0x5D, 0x0F, 0x3E, 0x0D, 0x3F, 0x03, 0x0E, 0x16, 0x34, 0x5F,
	0x00, 0x35, 0x21, 0x0E, 0x03, 0x22, 0x0E, 0x58, 0x36, 0x19, 0x3F, 0x77,
	0x3F, 0x22, 0x09, 0x28, 0x2D, 0x16, 0x0D, 0x1D, 0x3F, 0x0A, 0x03, 0x32,
	0x17, 0x28, 0x03, 0x3E, 0x25, 0x00, 0x28, 0x29, 0x02, 0x28, 0x1B, 0x23,
	0x21, 0x06, 0x02, 0x45, 0x07, 0x7A, 0x0A, 0x31, 0x3A, 0x27, 0x23, 0x5C,
	0x30, 0x05, 0x53, 0x75, 0x5E, 0x20, 0x5E, 0x53, 0x04, 0x0D, 0x03, 0x16,
	0x5F, 0x3B, 0x29, 0x05, 0x22, 0x0A, 0x73, 0x3D, 0x04, 0x09, 0x5A, 0x30,
	0x0D, 0x18, 0x57, 0x5D, 0x0F, 0x2F, 0x0C, 0x06, 0x32, 0x20, 0x0F, 0x0C,
	0x1B, 0x39, 0x29, 0x5E, 0x4E, 0x3F, 0x29, 0x0B, 0x14, 0x20, 0x58, 0x31,
	0x73, 0x5C, 0x52, 0x3B, 0x2E, 0x01, 0x5F, 0x51, 0x5D, 0x58, 0x1A, 0x5A,
	0x39, 0x41, 0x0D, 0x76, 0x5B, 0x0F, 0x27, 0x31, 0x1B, 0x26, 0x04, 0x0F,
	0x06, 0x3A, 0x1F, 0x31, 0x07, 0x39, 0x2E, 0x3C, 0x58, 0x26, 0x24, 0x10,
	0x03, 0x17, 0x3B, 0x2A, 0x05, 0x59, 0x2E, 0x1A, 0x0C, 0x72, 0x0B, 0x25,
	0x06, 0x3D, 0x18, 0x01, 0x2B, 0x1D, 0x3A, 0x77, 0x07, 0x3B, 0x3C, 0x3F,
	0x2B, 0x00, 0x24, 0x03, 0x26, 0x77, 0x21, 0x30, 0x2A, 0x5F, 0x11, 0x03,
	0x57, 0x23, 0x22, 0x00, 0x2F, 0x14, 0x03, 0x0C, 0x05, 0x27, 0x05, 0x3F,
	0x5E, 0x01, 0x47, 0x29, 0x25, 0x08, 0x03, 0x2B, 0x20, 0x25, 0x22, 0x15,
	0x25, 0x04, 0x36, 0x07, 0x03, 0x29, 0x2A, 0x2F, 0x08, 0x34, 0x5B, 0x05,
	0x04, 0x13, 0x16, 0x55, 0x1B, 0x59, 0x20, 0x28, 0x27, 0x57, 0x25, 0x40,
	0x01, 0x34, 0x08, 0x36, 0x2C, 0x0C, 0x0D, 0x16, 0x29, 0x25, 0x25, 0x09,
	0x50, 0x1A, 0x58, 0x0E, 0x47, 0x06, 0x3B, 0x23, 0x15, 0x5D, 0x10, 0x09,
	0x2E, 0x0D, 0x2E, 0x23, 0x20, 0x06, 0x00, 0x3F, 0x34, 0x2C, 0x2E, 0x2B,
	0x0B, 0x59, 0x29, 0x2F, 0x00, 0x5F, 0x12, 0x28, 0x02, 0x07, 0x28, 0x05,
	0x2B, 0x29, 0x24, 0x43, 0x27, 0x19, 0x58, 0x14, 0x1C, 0x3B, 0x3B, 0x3A,
	0x1A, 0x1B, 0x23, 0x5F, 0x20, 0x2E, 0x5B, 0x28, 0x07, 0x12, 0x24, 0x0A,
	0x20, 0x5E, 0x11, 0x03, 0x59, 0x07, 0x2D, 0x03, 0x75, 0x1F, 0x11, 0x20,
	0x2D, 0x74, 0x3E, 0x23, 0x34, 0x2F, 0x32, 0x00, 0x22, 0x2B, 0x19, 0x12,
	0x59, 0x17, 0x20, 0x38, 0x03, 0x08, 0x4E, 0x25, 0x26, 0x35, 0x0B, 0x08,
	0x1B, 0x03, 0x75, 0x05, 0x24, 0x01, 0x03, 0x05, 0x1E, 0x10, 0x27, 0x40,
	0x2C, 0x08, 0x56, 0x1C, 0x1B, 0x76, 0x24, 0x54, 0x2F, 0x32, 0x17, 0x1C,
	0x0A, 0x19, 0x24, 0x74, 0x0D, 0x2A, 0x08, 0x08, 0x24, 0x06, 0x34, 0x2F,
	0x44, 0x29, 0x20, 0x17, 0x2D, 0x5B, 0x23, 0x06, 0x07, 0x3A, 0x40, 0x25,
	0x18, 0x22, 0x04, 0x5B, 0x34, 0x05, 0x30, 0x0B, 0x2D, 0x3A, 0x3D, 0x11,
	0x5A, 0x02, 0x06, 0x3A, 0x56, 0x02, 0x44, 0x7A, 0x5C, 0x14, 0x5E, 0x52,
	0x08, 0x18, 0x28, 0x29, 0x38, 0x08, 0x2B, 0x36, 0x3A, 0x2A, 0x7B, 0x23,
	0x58, 0x59, 0x3E, 0x00, 0x21, 0x09, 0x1E, 0x59, 0x04, 0x26, 0x09, 0x0C,
	0x38, 0x00, 0x3F, 0x2D, 0x2C, 0x0D, 0x03, 0x06, 0x24, 0x00, 0x0E, 0x0B,
	0x0F, 0x35, 0x01, 0x5C, 0x2E, 0x36, 0x52, 0x21, 0x44, 0x1A, 0x34, 0x4A,
	0x34, 0x27, 0x7A, 0x01, 0x33, 0x2F, 0x32, 0x32, 0x0E, 0x3B, 0x29, 0x0A,
	0x10, 0x59, 0x32, 0x22, 0x07, 0x12, 0x27, 0x09, 0x57, 0x2C, 0x35, 0x3E,
	0x30, 0x3A, 0x5F, 0x0D, 0x0D, 0x2A, 0x5B, 0x53, 0x0B, 0x0A, 0x33, 0x1F,
	0x32, 0x05, 0x29, 0x06, 0x2A, 0x19, 0x0B, 0x26, 0x57, 0x22, 0x1E, 0x26,
	0x54, 0x09, 0x2C, 0x32, 0x09, 0x26, 0x0E, 0x2A, 0x5B, 0x0B, 0x07, 0x06,
	0x2A, 0x5D, 0x13, 0x02, 0x29, 0x20, 0x1F, 0x07, 0x5F, 0x20, 0x19, 0x1E,
	0x0E, 0x59, 0x05, 0x22, 0x1B, 0x2B, 0x0A, 0x27, 0x2C, 0x2C, 0x03, 0x2A,
	0x28, 0x2F, 0x58, 0x2A, 0x47, 0x24, 0x08, 0x20, 0x16, 0x3D, 0x59, 0x5E,
	0x5E, 0x2B, 0x2A, 0x58, 0x26, 0x28, 0x30, 0x01, 0x2D, 0x27, 0x09, 0x12,
	0x27, 0x25, 0x27, 0x44, 0x04, 0x1C, 0x0C, 0x21, 0x3F, 0x3A, 0x08, 0x0A,
	0x1D, 0x3D, 0x0A, 0x04, 0x54, 0x2D, 0x1F, 0x03, 0x0B, 0x2A, 0x20, 0x13,
	0x00, 0x35, 0x55, 0x58, 0x02, 0x2C, 0x0D, 0x24, 0x2B, 0x1F, 0x17, 0x3C,
	0x57, 0x25, 0x39, 0x03, 0x03, 0x59, 0x1B, 0x26, 0x0B, 0x2A, 0x13, 0x24,
	0x03, 0x77, 0x1F, 0x02, 0x05, 0x31, 0x71, 0x23, 0x58, 0x37, 0x25, 0x32,
	0x35, 0x32, 0x28, 0x03, 0x76, 0x39, 0x24, 0x06, 0x00, 0x24, 0x24, 0x33,
	0x04, 0x23, 0x06, 0x0A, 0x34, 0x2A, 0x28, 0x14, 0x05, 0x28, 0x04, 0x5B,
	0x2B, 0x35, 0x1B, 0x01, 0x02, 0x04, 0x35, 0x24, 0x41, 0x0A, 0x0D, 0x2F,
	0x16, 0x45, 0x27, 0x06, 0x2B, 0x38, 0x28, 0x39, 0x0E, 0x26, 0x58, 0x19,
	0x3D, 0x2B, 0x15, 0x2C, 0x2D, 0x3A, 0x25, 0x27, 0x59, 0x3D, 0x08, 0x13,
	0x25, 0x16, 0x3E, 0x3A, 0x0A, 0x47, 0x4E, 0x3E, 0x32, 0x12, 0x02, 0x24,
	0x16, 0x0C, 0x27, 0x29, 0x2C, 0x57, 0x2F, 0x29, 0x14, 0x28, 0x08, 0x2D,
	0x2B, 0x0B, 0x07, 0x34, 0x26, 0x0F, 0x27, 0x25, 0x3F, 0x18, 0x12, 0x06,
	0x16, 0x5E, 0x20, 0x10, 0x00, 0x59, 0x09, 0x1E, 0x04, 0x2B, 0x30, 0x21,
	0x1B, 0x2A, 0x47, 0x2A, 0x09, 0x1F, 0x03, 0x03, 0x18, 0x03, 0x3A, 0x07,
	0x2E, 0x35, 0x27, 0x01, 0x1B, 0x3B, 0x33, 0x27, 0x0A, 0x0E, 0x1B, 0x17,
	0x2D, 0x5B, 0x11, 0x14, 0x06, 0x07, 0x22, 0x2B, 0x58, 0x53, 0x20, 0x53,
	0x35, 0x07, 0x2E, 0x2D, 0x3A, 0x25, 0x26, 0x09, 0x08, 0x2C, 0x11, 0x58,
	0x0B, 0x16, 0x44, 0x28, 0x5F, 0x4A, 0x5D, 0x23, 0x18, 0x15, 0x05, 0x2C,
	0x2A, 0x31, 0x22, 0x19, 0x03, 0x53, 0x0D, 0x2A, 0x13, 0x3F, 0x5B, 0x29,
	0x39, 0x50, 0x2F, 0x1A, 0x2E, 0x58, 0x07, 0x29, 0x20, 0x6D, 0x00, 0x13,
	0x0A, 0x2F, 0x01, 0x0E, 0x24, 0x36, 0x2E, 0x13, 0x35, 0x02, 0x20, 0x53,
	0x76, 0x20, 0x30, 0x1E, 0x26, 0x2B, 0x0B, 0x38, 0x41, 0x3B, 0x0F, 0x26,
	0x23, 0x57, 0x26, 0x2C, 0x3A, 0x20, 0x08, 0x2A, 0x0D, 0x2E, 0x25, 0x14,
	0x5B, 0x14, 0x2B, 0x2C, 0x2B, 0x2F, 0x7B, 0x39, 0x33, 0x3C, 0x31, 0x7A,
	0x2E, 0x08, 0x1D, 0x39, 0x74, 0x03, 0x04, 0x3F, 0x22, 0x0D, 0x03, 0x32,
	0x59, 0x08, 0x12, 0x5A, 0x15, 0x14, 0x11, 0x75, 0x0E, 0x37, 0x25, 0x2A,
	0x17, 0x29, 0x55, 0x58, 0x05, 0x7A, 0x09, 0x27, 0x3D, 0x02, 0x30, 0x2D,
	0x06, 0x24, 0x40, 0x0D, 0x01, 0x25, 0x29, 0x25, 0x0E, 0x39, 0x23, 0x1F,
	0x2F, 0x07, 0x27, 0x11, 0x2F, 0x5A, 0x27, 0x29, 0x29, 0x2D, 0x39, 0x27,
	0x0A, 0x24, 0x3F, 0x32, 0x35, 0x28, 0x0B, 0x0B, 0x3B, 0x3B, 0x0B, 0x57,
	0x25, 0x28, 0x0B, 0x5C, 0x4E, 0x2B, 0x44, 0x74, 0x21, 0x0F, 0x09, 0x29,
	0x2B, 0x25, 0x27, 0x5A, 0x09, 0x2C, 0x03, 0x0C, 0x01, 0x38, 0x21, 0x14,
	0x30, 0x00, 0x13, 0x7A, 0x3B, 0x30, 0x16, 0x3A, 0x34, 0x2A, 0x59, 0x5A,
	0x22, 0x77, 0x0B, 0x33, 0x2B, 0x04, 0x2F, 0x3D, 0x56, 0x0D, 0x1C, 0x12,
	0x07, 0x22, 0x3C, 0x31, 0x70, 0x0D, 0x32, 0x2F, 0x11, 0x2B, 0x24, 0x0A,
	0x20, 0x0A, 0x2E, 0x18, 0x20, 0x34, 0x59, 0x0F, 0x02, 0x06, 0x58, 0x5C,
	0x0C, 0x39, 0x30, 0x39, 0x38, 0x17, 0x38, 0x20, 0x5A, 0x3E, 0x03, 0x15,
	0x24, 0x36, 0x25, 0x21, 0x3F, 0x2F, 0x5E, 0x18, 0x0F, 0x20, 0x18, 0x02,
	0x0C, 0x35, 0x3F, 0x16, 0x39, 0x11, 0x00, 0x55, 0x36, 0x0F, 0x26, 0x2B,
	0x0B, 0x12, 0x37, 0x12, 0x31, 0x2F, 0x08, 0x05, 0x2F, 0x2C, 0x09, 0x3B,
	0x0F, 0x3D, 0x32, 0x0D, 0x18, 0x3A, 0x1F, 0x03, 0x23, 0x22, 0x0D, 0x09,
	0x38, 0x24, 0x2C, 0x09, 0x06, 0x72, 0x27, 0x37, 0x06, 0x39, 0x75, 0x2A,
	0x35, 0x3F, 0x3B, 0x3B, 0x2B, 0x25, 0x3F, 0x3A, 0x2F, 0x3C, 0x2F, 0x17,
	0x18, 0x2F, 0x29, 0x33, 0x2F, 0x0E, 0x2F, 0x36, 0x06, 0x29, 0x08, 0x75,
	0x5A, 0x34, 0x29, 0x44, 0x30, 0x05, 0x04, 0x0F, 0x27, 0x11, 0x2A, 0x27,
	0x29, 0x5A, 0x17, 0x16, 0x2A, 0x2D, 0x3A, 0x2D, 0x21, 0x12, 0x07, 0x23,
	0x00, 0x3A, 0x0B, 0x29, 0x21, 0x3B, 0x1B, 0x04, 0x37, 0x0D, 0x07, 0x20,
	0x4E, 0x3C, 0x40, 0x0D, 0x1D, 0x38, 0x3F, 0x1A, 0x29, 0x39, 0x0D, 0x21,
	0x22, 0x15, 0x2D, 0x58, 0x22, 0x2A, 0x10, 0x2D, 0x25, 0x5E, 0x1E, 0x1A,
	0x0F, 0x51, 0x0B, 0x5D, 0x29, 0x26, 0x09, 0x23, 0x29, 0x34, 0x19, 0x2C,
	0x2D, 0x3A, 0x33, 0x23, 0x22, 0x18, 0x5E, 0x1A, 0x04, 0x15, 0x5D, 0x11,
	0x3B, 0x5E, 0x2D, 0x00, 0x1B, 0x15, 0x09, 0x2B, 0x1D, 0x1D, 0x74, 0x0F,
	0x29, 0x45, 0x11, 0x71, 0x0E, 0x2E, 0x5A, 0x0C, 0x0B, 0x3E, 0x30, 0x26,
	0x0D, 0x09, 0x06, 0x04, 0x0B, 0x1B, 0x01, 0x54, 0x18, 0x3C, 0x24, 0x2E,
	0x1C, 0x11, 0x29, 0x5A, 0x0B, 0x01, 0x17, 0x0D, 0x04, 0x18, 0x21, 0x13,
	0x5B, 0x19, 0x74, 0x08, 0x00, 0x05, 0x5A, 0x09, 0x2A, 0x07, 0x00, 0x5D,
	0x00, 0x2F, 0x09, 0x2F, 0x33, 0x29, 0x43, 0x27, 0x3E, 0x22, 0x70, 0x26,
	0x57, 0x3E, 0x06, 0x75, 0x2D, 0x07, 0x00, 0x33, 0x3B, 0x39, 0x09, 0x57,
	0x0C, 0x3A, 0x2E, 0x55, 0x07, 0x3D, 0x03, 0x3C, 0x30, 0x0F, 0x18, 0x00,
	0x24, 0x04, 0x1D, 0x01, 0x15, 0x0A, 0x0F, 0x16, 0x1B, 0x0B, 0x28, 0x08,
	0x1D, 0x19, 0x2F, 0x35, 0x05, 0x3A, 0x04, 0x71, 0x2E, 0x33, 0x1D, 0x28,
	0x6D, 0x5D, 0x0F, 0x0C, 0x08, 0x1B, 0x0E, 0x38, 0x5C, 0x3C, 0x0A, 0x29,
	0x07, 0x41, 0x39, 0x06, 0x07, 0x1B, 0x29, 0x09, 0x14, 0x25, 0x56, 0x3F,
	0x2A, 0x69, 0x3F, 0x33, 0x14, 0x26, 0x2C, 0x1E, 0x28, 0x04, 0x3F, 0x32,
	0x00, 0x14, 0x02, 0x5B, 0x16, 0x5C, 0x59, 0x58, 0x25, 0x32, 0x38, 0x2E,
	0x1A, 0x18, 0x2C, 0x07, 0x02, 0x24, 0x23, 0x24, 0x2F, 0x13, 0x3E, 0x2F,
	0x01, 0x2A, 0x51, 0x01, 0x05, 0x31, 0x1F, 0x35, 0x24, 0x27, 0x05, 0x59,
	0x0D, 0x1E, 0x03, 0x14, 0x26, 0x51, 0x39, 0x03, 0x71, 0x04, 0x09, 0x2A,
	0x5D, 0x73, 0x06, 0x18, 0x41, 0x31, 0x20, 0x15, 0x39, 0x5E, 0x21, 0x6D,
	0x1E, 0x2C, 0x18, 0x5D, 0x14, 0x1D, 0x37, 0x14, 0x39, 0x3A, 0x04, 0x22,
	0x2F, 0x13, 0x0B, 0x0D, 0x0A, 0x0C, 0x2A, 0x34, 0x2F, 0x05, 0x38, 0x22,
	0x70, 0x25, 0x14, 0x2B, 0x3D, 0x00, 0x26, 0x57, 0x05, 0x40, 0x6D, 0x27,
	0x55, 0x38, 0x1F, 0x3B, 0x43, 0x37, 0x2F, 0x24, 0x09, 0x3B, 0x30, 0x58,
	0x31, 0x10, 0x27, 0x10, 0x05, 0x25, 0x01, 0x0F, 0x09, 0x24, 0x1B, 0x1B,
	0x14, 0x50, 0x5B, 0x0E, 0x74, 0x24, 0x32, 0x19, 0x19, 0x28, 0x18, 0x23,
	0x2C, 0x3E, 0x0E, 0x35, 0x36, 0x04, 0x0A, 0x21, 0x3F, 0x3B, 0x34, 0x3C,
	0x2D, 0x3C, 0x29, 0x3A, 0x26, 0x69, 0x00, 0x24, 0x2C, 0x2E, 0x23, 0x03,
	0x08, 0x27, 0x1A, 0x18, 0x28, 0x57, 0x09, 0x53, 0x08, 0x0B, 0x25, 0x23,
	0x2A, 0x38, 0x06, 0x34, 0x5D, 0x1F, 0x76, 0x28, 0x33, 0x25, 0x3E, 0x33,
	0x47, 0x09, 0x5A, 0x0C, 0x2B, 0x00, 0x18, 0x34, 0x29, 0x06, 0x47, 0x51,
	0x5C, 0x29, 0x07, 0x3C, 0x0D, 0x3D, 0x2A, 0x2A, 0x07, 0x29, 0x0F, 0x08,
	0x27, 0x29, 0x27, 0x29, 0x0E, 0x28, 0x35, 0x30, 0x5A, 0x5D, 0x2C, 0x14,
	0x34, 0x2F, 0x00, 0x29, 0x59, 0x0C, 0x5F, 0x1C, 0x7B, 0x3D, 0x0F, 0x03,
	0x1A, 0x69, 0x06, 0x22, 0x05, 0x20, 0x0E, 0x26, 0x31, 0x2C, 0x2E, 0x17,
	0x23, 0x22, 0x3F, 0x5D, 0x17, 0x27, 0x12, 0x2C, 0x12, 0x2F, 0x25, 0x18,
	0x3C, 0x5F, 0x25, 0x39, 0x2B, 0x0D, 0x28, 0x06, 0x21, 0x07, 0x00, 0x03,
	0x25, 0x28, 0x31, 0x2D, 0x3A, 0x35, 0x27, 0x23, 0x1C, 0x18, 0x32, 0x26,
	0x27, 0x1A, 0x2A, 0x26, 0x5A, 0x28, 0x5A, 0x24, 0x73, 0x00, 0x20, 0x3F,
	0x02, 0x0E, 0x0B, 0x30, 0x22, 0x5D, 0x13, 0x00, 0x22, 0x14, 0x06, 0x32,
	0x0F, 0x31, 0x01, 0x29, 0x18, 0x2E, 0x03, 0x01, 0x1C, 0x35, 0x2E, 0x29,
	0x3A, 0x19, 0x0B, 0x22, 0x0D, 0x1E, 0x20, 0x27, 0x2E, 0x52, 0x3B, 0x5B,
	0x0C, 0x2E, 0x39, 0x41, 0x31, 0x21, 0x3C, 0x25, 0x21, 0x2A, 0x6D, 0x35,
	0x58, 0x25, 0x2F, 0x2A, 0x2D, 0x00, 0x3C, 0x38, 0x2E, 0x38, 0x24, 0x25,
	0x39, 0x10, 0x22, 0x35, 0x01, 0x1A, 0x2A, 0x05, 0x28, 0x0A, 0x05, 0x36,
	0x1F, 0x0C, 0x22, 0x0C, 0x38, 0x19, 0x00, 0x5D, 0x12, 0x76, 0x0E, 0x1B,
	0x5C, 0x59, 0x1A, 0x2F, 0x13, 0x26, 0x31, 0x18, 0x3F, 0x37, 0x58, 0x5C,
	0x75, 0x2E, 0x11, 0x19, 0x31, 0x34, 0x00, 0x24, 0x0B, 0x28, 0x23, 0x2D,
	0x12, 0x3A, 0x05, 0x36, 0x1F, 0x14, 0x19, 0x08, 0x0B, 0x0B, 0x1B, 0x0A,
	0x31, 0x26, 0x26, 0x17, 0x02, 0x25, 0x31, 0x19, 0x36, 0x19, 0x58, 0x21,
	0x1B, 0x05, 0x17, 0x24, 0x18, 0x55, 0x58, 0x24, 0x1D, 0x38, 0x5B, 0x28,
	0x19, 0x58, 0x3A, 0x3F, 0x14, 0x5C, 0x1C, 0x10, 0x15, 0x31, 0x0D, 0x2C,
	0x21, 0x3C, 0x57, 0x2D, 0x01, 0x28, 0x3E, 0x18, 0x20, 0x5E, 0x0D, 0x21,
	0x14, 0x19, 0x2A, 0x25, 0x3C, 0x2E, 0x5F, 0x1E, 0x08, 0x2B, 0x18, 0x36,
	0x3C, 0x13, 0x24, 0x0F, 0x2D, 0x0F, 0x3A, 0x00, 0x28, 0x08, 0x23, 0x31,
	0x2F, 0x38, 0x2D, 0x2F, 0x10, 0x3C, 0x58, 0x45, 0x52, 0x73, 0x54, 0x2E,
	0x1E, 0x2F, 0x29, 0x27, 0x0F, 0x2C, 0x09, 0x03, 0x06, 0x36, 0x2C, 0x19,
	0x11, 0x58, 0x16, 0x45, 0x23, 0x0A, 0x3D, 0x4E, 0x1F, 0x1C, 0x74, 0x5E,
	0x37, 0x09, 0x0C, 0x7B, 0x19, 0x0A, 0x22, 0x1A, 0x25, 0x09, 0x57, 0x24,
	0x0F, 0x27, 0x54, 0x26, 0x3D, 0x32, 0x30, 0x34, 0x55, 0x0A, 0x1F, 0x08,
	0x34, 0x33, 0x41, 0x12, 0x07, 0x5B, 0x24, 0x3B, 0x3A, 0x12, 0x07, 0x2C,
	0x0B, 0x31, 0x77, 0x2D, 0x22, 0x3F, 0x3F, 0x23, 0x01, 0x35, 0x19, 0x2A,
	0x73, 0x15, 0x36, 0x3C, 0x1B, 0x07, 0x2E, 0x13, 0x0B, 0x5A, 0x2A, 0x27,
	0x54, 0x5D, 0x06, 0x09, 0x07, 0x22, 0x0A, 0x1C, 0x74, 0x21, 0x2A, 0x2D,
	0x5D, 0x0F, 0x0F, 0x35, 0x5C, 0x23, 0x13, 0x1F, 0x32, 0x09, 0x20, 0x15,
	0x29, 0x2D, 0x2C, 0x11, 0x13, 0x09, 0x12, 0x2D, 0x05, 0x10, 0x1F, 0x53,
	0x0D, 0x08, 0x21, 0x38, 0x38, 0x1D, 0x00, 0x38, 0x01, 0x16, 0x5D, 0x06,
	0x37, 0x5B, 0x0D, 0x1D, 0x1F, 0x0F, 0x3E, 0x23, 0x06, 0x58, 0x0F, 0x58,
	0x0B, 0x28, 0x39, 0x28, 0x21, 0x2C, 0x14, 0x24, 0x38, 0x18, 0x56, 0x21,
	0x1C, 0x21, 0x5B, 0x33, 0x14, 0x18, 0x2C, 0x23, 0x53, 0x0D, 0x5C, 0x04,
	0x16, 0x15, 0x36, 0x24, 0x38, 0x0F, 0x55, 0x0A, 0x39, 0x0C, 0x02, 0x03,
	0x21, 0x52, 0x25, 0x5B, 0x53, 0x04, 0x1D, 0x18, 0x23, 0x58, 0x1B, 0x5C,
	0x70, 0x20, 0x17, 0x0F, 0x1E, 0x7B, 0x01, 0x56, 0x09, 0x5B, 0x16, 0x5E,
	0x25, 0x09, 0x5F, 0x0D, 0x06, 0x06, 0x5B, 0x24, 0x06, 0x1F, 0x55, 0x21,
	0x27, 0x25, 0x5A, 0x14, 0x2A, 0x06, 0x76, 0x23, 0x56, 0x1B, 0x2A, 0x73,
	0x09, 0x51, 0x0D, 0x23, 0x10, 0x5C, 0x05, 0x26, 0x21, 0x72, 0x08, 0x0F,
	0x3C, 0x13, 0x26, 0x24, 0x37, 0x5E, 0x08, 0x71, 0x3E, 0x52, 0x0B, 0x3A,
	0x29, 0x0E, 0x53, 0x3A, 0x0C, 0x77, 0x23, 0x0B, 0x05, 0x5E, 0x0D, 0x38,
	0x12, 0x5B, 0x24, 0x0E, 0x07, 0x57, 0x1B, 0x3F, 0x2F, 0x59, 0x2C, 0x59,
	0x12, 0x0C, 0x1E, 0x04, 0x5C, 0x08, 0x0A, 0x36, 0x51, 0x0A, 0x05, 0x08,
	0x5E, 0x05, 0x00, 0x31, 0x3A, 0x08, 0x0F, 0x38, 0x59, 0x21, 0x5F, 0x3B,
	0x26, 0x39, 0x10, 0x01, 0x56, 0x45, 0x27, 0x25, 0x58, 0x14, 0x04, 0x02,
	0x77, 0x23, 0x2D, 0x1D, 0x5F, 0x37, 0x20, 0x08, 0x58, 0x1E, 0x0E, 0x01,
	0x55, 0x09, 0x5D, 0x09, 0x18, 0x52, 0x0A, 0x5A, 0x21, 0x24, 0x37, 0x5E,
	0x0F, 0x1A, 0x26, 0x50, 0x0A, 0x05, 0x14, 0x14, 0x05, 0x36, 0x3D, 0x73,
	0x0F, 0x52, 0x3B, 0x23, 0x01, 0x22, 0x0C, 0x59, 0x24, 0x20, 0x0B, 0x54,
	0x1B, 0x01, 0x2F, 0x59, 0x2E, 0x0C, 0x1E, 0x77, 0x19, 0x2D, 0x03, 0x5D,
	0x37, 0x0E, 0x0C, 0x5B, 0x2A, 0x3A, 0x38, 0x15, 0x5D, 0x39, 0x71, 0x0F,
	0x29, 0x0A, 0x59, 0x26, 0x5F, 0x2B, 0x5D, 0x0F, 0x1A, 0x08, 0x19, 0x0A,
	0x58, 0x26, 0x5F, 0x02, 0x5D, 0x0F, 0x71, 0x00, 0x4E, 0x0D, 0x11, 0x0D,
	0x5F, 0x12, 0x26, 0x39, 0x3B, 0x08, 0x0F, 0x28, 0x5A, 0x21, 0x5E, 0x05,
	0x00, 0x31, 0x2B, 0x39, 0x1B, 0x2B, 0x07, 0x08, 0x38, 0x34, 0x1B, 0x0D,
	0x2F, 0x26, 0x26, 0x34, 0x13, 0x27, 0x3A, 0x0D, 0x3A, 0x40, 0x0B, 0x20,
	0x09, 0x25, 0x20, 0x21, 0x5F, 0x2D, 0x14, 0x53, 0x3B, 0x3A, 0x09, 0x19,
	0x26, 0x0D, 0x0E, 0x17, 0x04, 0x44, 0x2C, 0x16, 0x12, 0x20, 0x03, 0x1B,
	0x38, 0x22, 0x2A, 0x2A, 0x0F, 0x06, 0x2A, 0x19, 0x00, 0x00, 0x2D, 0x12,
	0x25, 0x1C, 0x36, 0x20, 0x32, 0x56, 0x24, 0x1B, 0x38, 0x26, 0x14, 0x18,
	0x15, 0x2F, 0x16, 0x5B, 0x2C, 0x10, 0x1A, 0x2F, 0x19, 0x5B, 0x23, 0x3C,
	0x19, 0x00, 0x21, 0x77, 0x3B, 0x26, 0x5A, 0x1E, 0x11, 0x2D, 0x58, 0x08,
	0x53, 0x03, 0x08, 0x31, 0x5A, 0x20, 0x0C, 0x07, 0x26, 0x2B, 0x32, 0x10,
	0x43, 0x17, 0x2F, 0x0D, 0x06, 0x5C, 0x38, 0x02, 0x0C, 0x74, 0x14, 0x20,
	0x34, 0x18, 0x07, 0x54, 0x03, 0x04, 0x22, 0x75, 0x24, 0x55, 0x1D, 0x3E,
	0x21, 0x3D, 0x30, 0x3F, 0x13, 0x2C, 0x2F, 0x32, 0x1B, 0x32, 0x13, 0x1A,
	0x2C, 0x05, 0x58, 0x07, 0x3E, 0x54, 0x5A, 0x2A, 0x24, 0x06, 0x0E, 0x2B,
	0x2E, 0x15, 0x2E, 0x57, 0x17, 0x2E, 0x21, 0x09, 0x24, 0x36, 0x1B, 0x28,
	0x26, 0x2B, 0x1D, 0x19, 0x1B, 0x1A, 0x31, 0x2C, 0x32, 0x72, 0x58, 0x08,
	0x26, 0x58, 0x2C, 0x2D, 0x37, 0x2D, 0x53, 0x32, 0x28, 0x07, 0x23, 0x29,
	0x1B, 0x05, 0x2C, 0x3A, 0x40, 0x07, 0x29, 0x22, 0x23, 0x26, 0x17, 0x2F,
	0x4E, 0x14, 0x27, 0x38, 0x21, 0x33, 0x57, 0x39, 0x33, 0x07, 0x06, 0x09,
	0x13, 0x01, 0x25, 0x20, 0x27, 0x58, 0x09, 0x15, 0x24, 0x04, 0x07, 0x7A,
	0x20, 0x25, 0x3C, 0x21, 0x3B, 0x25, 0x2C, 0x19, 0x29, 0x0F, 0x15, 0x36,
	0x3B, 0x32, 0x13, 0x43, 0x2B, 0x5A, 0x05, 0x35, 0x14, 0x26, 0x29, 0x3A,
	0x11, 0x38, 0x22, 0x0C, 0x39, 0x0E, 0x35, 0x30, 0x1D, 0x5B, 0x2C, 0x27,
	0x32, 0x1D, 0x32, 0x0B, 0x01, 0x0F, 0x3A, 0x3A, 0x74, 0x24, 0x59, 0x09,
	0x44, 0x72, 0x08, 0x0F, 0x5B, 0x0A, 0x17, 0x00, 0x3B, 0x09, 0x00, 0x7A,
	0x1F, 0x03, 0x2B, 0x24, 0x2F, 0x34, 0x3B, 0x1D, 0x31, 0x2C, 0x3D, 0x57,
	0x25, 0x12, 0x31, 0x07, 0x2B, 0x14, 0x23, 0x01, 0x5F, 0x32, 0x56, 0x13,
	0x0F, 0x29, 0x25, 0x2B, 0x11, 0x30, 0x09, 0x07, 0x07, 0x22, 0x71, 0x23,
	0x18, 0x2B, 0x1E, 0x0E, 0x16, 0x23, 0x25, 0x24, 0x16, 0x20, 0x28, 0x3E,
	0x5E, 0x76, 0x34, 0x29, 0x04, 0x2A, 0x3A, 0x25, 0x12, 0x06, 0x44, 0x36,
	0x2F, 0x03, 0x03, 0x5F, 0x2F, 0x15, 0x32, 0x5F, 0x1C, 0x74, 0x16, 0x05,
	0x2F, 0x3E, 0x21, 0x59, 0x14, 0x09, 0x22, 0x69, 0x0F, 0x0F, 0x28, 0x11,
	0x26, 0x02, 0x28, 0x28, 0x01, 0x05, 0x24, 0x0F, 0x3C, 0x04, 0x3A, 0x38,
	0x30, 0x5A, 0x21, 0x01, 0x2D, 0x0E, 0x06, 0x03, 0x3B, 0x14, 0x13, 0x58,
	0x5F, 0x01, 0x2E, 0x26, 0x04, 0x2D, 0x2C, 0x15, 0x20, 0x0D, 0x1C, 0x05,
	0x47, 0x26, 0x19, 0x2A, 0x25, 0x28, 0x29, 0x01, 0x23, 0x77, 0x14, 0x55,
	0x23, 0x08, 0x0E, 0x28, 0x30, 0x56, 0x3B, 0x75, 0x2D, 0x30, 0x56, 0x08,
	0x0C, 0x5D, 0x57, 0x5C, 0x12, 0x74, 0x28, 0x2D, 0x0C, 0x06, 0x70, 0x34,
	0x26, 0x0C, 0x0F, 0x70, 0x3D, 0x26, 0x57, 0x1B, 0x37, 0x54, 0x1B, 0x1A,
	0x31, 0x13, 0x08, 0x34, 0x45, 0x5F, 0x0D, 0x0E, 0x23, 0x0A, 0x27, 0x12,
	0x47, 0x15, 0x3F, 0x1E, 0x72, 0x43, 0x54, 0x2D, 0x1C, 0x06, 0x54, 0x54,
	0x36, 0x3C, 0x15, 0x36, 0x03, 0x24, 0x5D, 0x11, 0x38, 0x2F, 0x0F, 0x26,
	0x3B, 0x5E, 0x33, 0x5D, 0x31, 0x0D, 0x5E, 0x18, 0x36, 0x24, 0x03, 0x19,
	0x15, 0x26, 0x08, 0x7A, 0x5B, 0x4E, 0x56, 0x31, 0x3B, 0x29, 0x0E, 0x2F,
	0x1A, 0x72, 0x02, 0x55, 0x24, 0x58, 0x24, 0x5D, 0x33, 0x59, 0x1D, 0x0F,
	0x2E, 0x13, 0x04, 0x08, 0x2C, 0x47, 0x53, 0x17, 0x02, 0x33, 0x43, 0x15,
	0x1D, 0x03, 0x12, 0x0A, 0x53, 0x03, 0x33, 0x75, 0x1A, 0x0F, 0x3F, 0x53,
	0x20, 0x1B, 0x35, 0x21, 0x11, 0x7A, 0x22, 0x36, 0x03, 0x21, 0x15, 0x22,
	0x53, 0x34, 0x22, 0x06, 0x5D, 0x32, 0x56, 0x0A, 0x06, 0x1B, 0x09, 0x1A,
	0x1E, 0x2B, 0x5C, 0x05, 0x07, 0x1C, 0x35, 0x23, 0x59, 0x19, 0x53, 0x09,
	0x14, 0x18, 0x27, 0x31, 0x35, 0x3B, 0x29, 0x3F, 0x01, 0x3B, 0x3A, 0x1B,
	0x5A, 0x2D, 0x2D, 0x59, 0x0F, 0x2A, 0x2E, 0x11, 0x35, 0x19, 0x3F, 0x5E,
	0x21, 0x24, 0x05, 0x2B, 0x2A, 0x38, 0x2B, 0x39, 0x14, 0x29, 0x23, 0x15,
	0x55, 0x39, 0x0C, 0x29, 0x3A, 0x2A, 0x16, 0x20, 0x03, 0x5A, 0x0F, 0x03,
	0x39, 0x21, 0x08, 0x18, 0x2B, 0x5B, 0x2E, 0x47, 0x24, 0x3F, 0x28, 0x2E,
	0x04, 0x20, 0x23, 0x5E, 0x2A, 0x1A, 0x0B, 0x2D, 0x0C, 0x0B, 0x25, 0x0A,
	0x2D, 0x1B, 0x1B, 0x08, 0x38, 0x59, 0x04, 0x11, 0x1D, 0x30, 0x0D, 0x04,
	0x29, 0x47, 0x2C, 0x5C, 0x44, 0x01, 0x3D, 0x2D, 0x0C, 0x5C, 0x0E, 0x3F,
	0x23, 0x09, 0x5F, 0x23, 0x1B, 0x0E, 0x37, 0x0D, 0x15, 0x47, 0x27, 0x34,
	0x0E, 0x71, 0x1A, 0x06, 0x5A, 0x2A, 0x07, 0x26, 0x2F, 0x00, 0x2F, 0x16,
	0x0B, 0x2A, 0x1B, 0x2C, 0x75, 0x58, 0x2C, 0x23, 0x1B, 0x25, 0x2B, 0x29,
	0x09, 0x5B, 0x3A, 0x1B, 0x0A, 0x2F, 0x00, 0x0D, 0x21, 0x12, 0x26, 0x29,
	0x0B, 0x25, 0x55, 0x2A, 0x03, 0x13, 0x28, 0x39, 0x2F, 0x00, 0x76, 0x34,
	0x2E, 0x29, 0x3B, 0x25, 0x5A, 0x2C, 0x2F, 0x29, 0x1A, 0x3D, 0x38, 0x26,
	0x02, 0x25, 0x2F, 0x04, 0x09, 0x3B, 0x71, 0x5E, 0x2B, 0x16, 0x44, 0x2C,
	0x00, 0x35, 0x1C, 0x03, 0x08, 0x0F, 0x05, 0x20, 0x01, 0x2A, 0x47, 0x37,
	0x5F, 0x29, 0x0C, 0x39, 0x32, 0x28, 0x13, 0x14, 0x3F, 0x07, 0x5F, 0x2F,
	0x28, 0x0F, 0x30, 0x0C, 0x24, 0x25, 0x5F, 0x32, 0x0F, 0x31, 0x08, 0x23,
	0x08, 0x5D, 0x3F, 0x23, 0x1C, 0x2B, 0x3E, 0x44, 0x0D, 0x18, 0x05, 0x0C,
	0x1B, 0x14, 0x22, 0x04, 0x58, 0x1B, 0x71, 0x09, 0x09, 0x45, 0x07, 0x32,
	0x26, 0x22, 0x5C, 0x0C, 0x6D, 0x0B, 0x2C, 0x41, 0x2C, 0x29, 0x21, 0x13,
	0x00, 0x44, 0x06, 0x06, 0x59, 0x19, 0x2F, 0x25, 0x58, 0x2F, 0x39, 0x1A,
	0x28, 0x1F, 0x20, 0x20, 0x2A, 0x7A, 0x58, 0x31, 0x21, 0x2C, 0x28, 0x2F,
	0x27, 0x5D, 0x5C, 0x0E, 0x0B, 0x2E, 0x18, 0x1A, 0x08, 0x0F, 0x23, 0x1A,
	0x2A, 0x0D, 0x58, 0x2C, 0x0D, 0x3B, 0x06, 0x03, 0x12, 0x0A, 0x27, 0x6D,
	0x14, 0x38, 0x45, 0x23, 0x27, 0x28, 0x04, 0x00, 0x5A, 0x0F, 0x5D, 0x33,
	0x1B, 0x01, 0x2C, 0x00, 0x03, 0x01, 0x5C, 0x23, 0x16, 0x39, 0x36, 0x44,
	0x74, 0x09, 0x13, 0x1E, 0x32, 0x70, 0x1D, 0x10, 0x58, 0x02, 0x2D, 0x0D,
	0x37, 0x2B, 0x5A, 0x2E, 0x20, 0x38, 0x1F, 0x59, 0x29, 0x0B, 0x54, 0x21,
	0x22, 0x7A, 0x1E, 0x27, 0x21, 0x44, 0x11, 0x15, 0x4E, 0x58, 0x44, 0x7A,
	0x1A, 0x28, 0x2F, 0x09, 0x13, 0x39, 0x2A, 0x5B, 0x23, 0x73, 0x5A, 0x59,
	0x59, 0x3A, 0x35, 0x0F, 0x17, 0x23, 0x3B, 0x0F, 0x2A, 0x35, 0x09, 0x58,
	0x76, 0x23, 0x20, 0x09, 0x29, 0x1B, 0x43, 0x2E, 0x19, 0x0D, 0x1B, 0x0F,
	0x25, 0x1E, 0x11, 0x2C, 0x0A, 0x54, 0x26, 0x58, 0x30, 0x43, 0x13, 0x3C,
	0x5C, 0x6D, 0x04, 0x2B, 0x14, 0x04, 0x26, 0x3D, 0x0D, 0x5A, 0x33, 0x17,
	0x04, 0x11, 0x1D, 0x09, 0x0B, 0x2B, 0x4E, 0x2C, 0x11, 0x13, 0x09, 0x30,
	0x18, 0x40, 0x03, 0x01, 0x23, 0x58, 0x03, 0x24, 0x1B, 0x51, 0x5E, 0x22,
	0x29, 0x22, 0x07, 0x09, 0x1B, 0x25, 0x0D, 0x35, 0x36, 0x5E, 0x10, 0x26,
	0x29, 0x00, 0x1B, 0x01, 0x23, 0x0B, 0x08, 0x00, 0x10, 0x43, 0x0B, 0x3C,
	0x23, 0x37, 0x1E, 0x0B, 0x0D, 0x3B, 0x0F, 0x28, 0x54, 0x2B, 0x5B, 0x74,
	0x3E, 0x17, 0x3C, 0x09, 0x23, 0x29, 0x24, 0x2C, 0x53, 0x2B, 0x02, 0x34,
	0x1F, 0x0A, 0x0A, 0x08, 0x0D, 0x37, 0x23, 0x03, 0x28, 0x30, 0x27, 0x24,
	0x2B, 0x0B, 0x22, 0x5A, 0x0A, 0x25, 0x02, 0x0D, 0x23, 0x24, 0x16, 0x04,
	0x0E, 0x0D, 0x2F, 0x00, 0x2F, 0x54, 0x1A, 0x1F, 0x25, 0x25, 0x2F, 0x59,
	0x24, 0x37, 0x28, 0x34, 0x2F, 0x44, 0x18, 0x59, 0x04, 0x2F, 0x09, 0x0E,
	0x54, 0x35, 0x08, 0x5A, 0x24, 0x07, 0x17, 0x21, 0x22, 0x71, 0x3E, 0x2F,
	0x2D, 0x2E, 0x25, 0x02, 0x0E, 0x3A, 0x08, 0x08, 0x01, 0x59, 0x00, 0x5E,
	0x10, 0x2E, 0x06, 0x34, 0x19, 0x2A, 0x14, 0x20, 0x19, 0x2A, 0x13, 0x15,
	0x0F, 0x2D, 0x59, 0x12, 0x26, 0x4A, 0x28, 0x0A, 0x07, 0x1C, 0x55, 0x03,
	0x32, 0x16, 0x5C, 0x2B, 0x5D, 0x5E, 0x0B, 0x3D, 0x37, 0x24, 0x32, 0x2D,
	0x04, 0x55, 0x3C, 0x59, 0x08, 0x2D, 0x1B, 0x1C, 0x5A, 0x1A, 0x34, 0x04,
	0x27, 0x1D, 0x6D, 0x3E, 0x36, 0x56, 0x05, 0x7A, 0x34, 0x54, 0x2C, 0x5F,
	0x11, 0x0F, 0x0F, 0x56, 0x38, 0x07, 0x0B, 0x0F, 0x5A, 0x52, 0x27, 0x5E,
	0x24, 0x26, 0x2A, 0x12, 0x2F, 0x36, 0x29, 0x09, 0x26, 0x23, 0x54, 0x5D,
	0x0C, 0x72, 0x05, 0x0E, 0x3D, 0x00, 0x08, 0x58, 0x50, 0x19, 0x20, 0x29,
	0x20, 0x56, 0x36, 0x09, 0x16, 0x5A, 0x52, 0x0C, 0x3F, 0x75, 0x5F, 0x03,
	0x3A, 0x5C, 0x1A, 0x0E, 0x25, 0x45, 0x27, 0x76, 0x29, 0x59, 0x17, 0x2F,
	0x34, 0x0B, 0x29, 0x5D, 0x29, 0x20, 0x06, 0x57, 0x0C, 0x04, 0x74, 0x0F,
	0x4E, 0x03, 0x2D, 0x3B, 0x09, 0x23, 0x18, 0x2E, 0x26, 0x34, 0x03, 0x39,
	0x31, 0x0E, 0x1B, 0x02, 0x17, 0x1E, 0x26, 0x3C, 0x59, 0x18, 0x07, 0x1B,
	0x28, 0x57, 0x14, 0x19, 0x34, 0x29, 0x0A, 0x45, 0x27, 0x76, 0x21, 0x4E,
	0x17, 0x20, 0x7B, 0x0D, 0x3B, 0x24, 0x0C, 0x2F, 0x06, 0x59, 0x08, 0x5C,
	0x09, 0x3C, 0x39, 0x38, 0x26, 0x23, 0x0D, 0x38, 0x57, 0x01, 0x01, 0x07,
	0x0C, 0x0B, 0x0C, 0x32, 0x1D, 0x54, 0x00, 0x5A, 0x73, 0x19, 0x54, 0x1E,
	0x31, 0x09, 0x2F, 0x13, 0x5C, 0x00, 0x36, 0x20, 0x39, 0x5E, 0x3C, 0x16,
	0x1D, 0x10, 0x29, 0x24, 0x23, 0x22, 0x10, 0x34, 0x1C, 0x0E, 0x05, 0x03,
	0x05, 0x19, 0x36, 0x55, 0x29, 0x5A, 0x1A, 0x2C, 0x14, 0x53, 0x2D, 0x23,
	0x25, 0x34, 0x52, 0x5F, 0x07, 0x0E, 0x5D, 0x12, 0x06, 0x5E, 0x2E, 0x0E,
	0x25, 0x5D, 0x23, 0x31, 0x58, 0x35, 0x17, 0x04, 0x2C, 0x5A, 0x0C, 0x16,
	0x1D, 0x2A, 0x36, 0x50, 0x06, 0x20, 0x36, 0x08, 0x56, 0x45, 0x2D, 0x15,
	0x2A, 0x13, 0x01, 0x59, 0x03, 0x58, 0x38, 0x0F, 0x24, 0x26, 0x2A, 0x56,
	0x0F, 0x19, 0x30, 0x5C, 0x12, 0x1F, 0x3F, 0x73, 0x22, 0x1B, 0x3A, 0x3F,
	0x0F, 0x22, 0x24, 0x16, 0x3E, 0x0C, 0x08, 0x36, 0x3B, 0x5F, 0x1A, 0x03,
	0x2A, 0x1B, 0x0A, 0x05, 0x2B, 0x2C, 0x27, 0x09, 0x00, 0x5F, 0x0B, 0x06,
	0x2C, 0x0B, 0x3B, 0x24, 0x17, 0x1F, 0x71, 0x2F, 0x50, 0x29, 0x5E, 0x2A,
	0x00, 0x36, 0x5B, 0x03, 0x73, 0x3B, 0x54, 0x06, 0x22, 0x0F, 0x05, 0x34,
	0x0D, 0x28, 0x17, 0x00, 0x22, 0x00, 0x39, 0x09, 0x2A, 0x28, 0x1F, 0x12,
	0x0A, 0x29, 0x2B, 0x26, 0x3E, 0x14, 0x0D, 0x0C, 0x17, 0x02, 0x04, 0x5C,
	0x18, 0x02, 0x38, 0x33, 0x05, 0x09, 0x16, 0x28, 0x10, 0x5D, 0x37, 0x3C,
	0x3E, 0x18, 0x3A, 0x25, 0x58, 0x2D, 0x10, 0x39, 0x37, 0x0A, 0x3C, 0x35,
	0x35, 0x14, 0x41, 0x3F, 0x7B, 0x20, 0x34, 0x24, 0x11, 0x20, 0x1D, 0x37,
	0x37, 0x0D, 0x14, 0x5E, 0x04, 0x59, 0x27, 0x24, 0x1D, 0x12, 0x5F, 0x02,
	0x73, 0x00, 0x0D, 0x1B, 0x38, 0x18, 0x21, 0x00, 0x22, 0x13, 0x71, 0x38,
	0x54, 0x28, 0x0A, 0x14, 0x5D, 0x57, 0x34, 0x08, 0x74, 0x02, 0x4E, 0x39,
	0x44, 0x09, 0x43, 0x0A, 0x1E, 0x5F, 0x1B, 0x20, 0x28, 0x5C, 0x53, 0x76,
	0x24, 0x33, 0x2C, 0x40, 0x73, 0x26, 0x13, 0x2A, 0x1E, 0x28, 0x14, 0x51,
	0x3C, 0x40, 0x23, 0x1E, 0x31, 0x07, 0x1D, 0x28, 0x5B, 0x06, 0x5E, 0x44,
	0x1A, 0x1A, 0x23, 0x2A, 0x0A, 0x20, 0x1C, 0x17, 0x3A, 0x0D, 0x6D, 0x5D,
	0x08, 0x37, 0x44, 0x73, 0x59, 0x55, 0x0D, 0x58, 0x0D, 0x23, 0x1B, 0x04,
	0x1D, 0x7B, 0x09, 0x38, 0x3E, 0x0D, 0x0E, 0x05, 0x55, 0x29, 0x5B, 0x16,
	0x34, 0x4E, 0x34, 0x0A, 0x12, 0x1A, 0x00, 0x21, 0x13, 0x7B, 0x24, 0x2B,
	0x5D, 0x5A, 0x10, 0x01, 0x23, 0x24, 0x1C, 0x24, 0x19, 0x22, 0x00, 0x07,
	0x27, 0x35, 0x4E, 0x28, 0x5B, 0x1B, 0x5C, 0x14, 0x06, 0x58, 0x0B, 0x47,
	0x57, 0x5F, 0x38, 0x07, 0x34, 0x2D, 0x26, 0x31, 0x3A, 0x34, 0x50, 0x1A,
	0x1E, 0x2C, 0x1E, 0x22, 0x2F, 0x5D, 0x69, 0x38, 0x33, 0x0B, 0x58, 0x76,
	0x22, 0x2B, 0x41, 0x1A, 0x24, 0x19, 0x17, 0x37, 0x01, 0x6D, 0x38, 0x0C,
	0x04, 0x09, 0x77, 0x01, 0x17, 0x5D, 0x0D, 0x11, 0x23, 0x52, 0x38, 0x13,
	0x72, 0x2D, 0x36, 0x1C, 0x19, 0x27, 0x07, 0x15, 0x24, 0x18, 0x36, 0x05,
	0x03, 0x59, 0x18, 0x24, 0x15, 0x07, 0x57, 0x20, 0x0E, 0x3B, 0x2E, 0x0D,
	0x18, 0x7B, 0x06, 0x28, 0x0B, 0x3C, 0x23, 0x5C, 0x2A, 0x21, 0x1A, 0x2F,
	0x54, 0x51, 0x26, 0x39, 0x08, 0x47, 0x52, 0x17, 0x5F, 0x0E, 0x47, 0x15,
	0x0A, 0x59, 0x20, 0x55, 0x51, 0x5D, 0x0D, 0x14, 0x47, 0x31, 0x1B, 0x0E,
	0x08, 0x1B, 0x11, 0x41, 0x3E, 0x29, 0x1E, 0x59, 0x14, 0x0C, 0x38, 0x35,
	0x0A, 0x3E, 0x3F, 0x07, 0x35, 0x24, 0x26, 0x2E, 0x26, 0x0F, 0x07, 0x57,
	0x0C, 0x25, 0x47, 0x00, 0x05, 0x07, 0x05, 0x34, 0x09, 0x03, 0x11, 0x12,
	0x0D, 0x2E, 0x5C, 0x52, 0x1B, 0x18, 0x1B, 0x0A, 0x32, 0x21, 0x09, 0x0C,
	0x08, 0x2D, 0x27, 0x08, 0x26, 0x38, 0x0C, 0x75, 0x0D, 0x29, 0x3E, 0x1A,
	0x2B, 0x59, 0x54, 0x22, 0x32, 0x2F, 0x5A, 0x54, 0x26, 0x18, 0x75, 0x55,
	0x30, 0x1E, 0x18, 0x20, 0x09, 0x15, 0x38, 0x59, 0x0C, 0x47, 0x4A, 0x20,
	0x59, 0x18, 0x1E, 0x55, 0x06, 0x12, 0x0C, 0x23, 0x35, 0x34, 0x3D, 0x2A,
	0x07, 0x28, 0x2A, 0x0C, 0x32, 0x5C, 0x1B, 0x45, 0x3D, 0x0E, 0x1E, 0x58,
	0x2D, 0x21, 0x75, 0x2D, 0x12, 0x2A, 0x1A, 0x31, 0x5A, 0x1B, 0x16, 0x0E,
	0x35, 0x3F, 0x55, 0x37, 0x22, 0x13, 0x09, 0x09, 0x22, 0x02, 0x0F, 0x2A,
	0x16, 0x02, 0x21, 0x71, 0x29, 0x29, 0x2B, 0x2C, 0x73, 0x22, 0x14, 0x36,
	0x03, 0x2A, 0x39, 0x17, 0x36, 0x04, 0x32, 0x04, 0x0B, 0x14, 0x5E, 0x10,
	0x1F, 0x38, 0x18, 0x27, 0x2A, 0x5E, 0x27, 0x3E, 0x25, 0x11, 0x3C, 0x09,
	0x2C, 0x02, 0x70, 0x21, 0x54, 0x20, 0x23, 0x0D, 0x5B, 0x53, 0x20, 0x32,
	0x3A, 0x5B, 0x0F, 0x04, 0x31, 0x00, 0x26, 0x2A, 0x17, 0x32, 0x17, 0x21,
	0x0C, 0x2C, 0x44, 0x7A, 0x15, 0x02, 0x45, 0x3D, 0x35, 0x02, 0x1B, 0x06,
	0x2F, 0x69, 0x39, 0x2F, 0x08, 0x11, 0x00, 0x43, 0x4A, 0x27, 0x25, 0x2E,
	0x1B, 0x23, 0x56, 0x04, 0x00, 0x47, 0x50, 0x3C, 0x00, 0x2F, 0x54, 0x26,
	0x5E, 0x52, 0x73, 0x58, 0x20, 0x5F, 0x58, 0x24, 0x19, 0x2B, 0x37, 0x0D,
	0x1B, 0x0B, 0x18, 0x5B, 0x58, 0x1A, 0x19, 0x18, 0x59, 0x04, 0x27, 0x14,
	0x2C, 0x27, 0x3B, 0x38, 0x0A, 0x19, 0x39, 0x3D, 0x35, 0x5C, 0x2A, 0x1F,
	0x0E, 0x27, 0x55, 0x0F, 0x3F, 0x2C, 0x29, 0x5A, 0x04, 0x5D, 0x1C, 0x27,
	0x25, 0x16, 0x05, 0x3E, 0x29, 0x1E, 0x19, 0x5B, 0x44, 0x74, 0x2A, 0x0C,
	0x27, 0x26, 0x74, 0x00, 0x38, 0x1B, 0x3E, 0x00, 0x18, 0x03, 0x3E, 0x03,
	0x33, 0x43, 0x2B, 0x20, 0x0A, 0x2A, 0x5E, 0x4E, 0x34, 0x1D, 0x08, 0x54,
	0x16, 0x5F, 0x09, 0x3B, 0x0A, 0x28, 0x21, 0x3A, 0x12, 0x22, 0x4E, 0x09,
	0x3F, 0x18, 0x59, 0x17, 0x5E, 0x28, 0x06, 0x3C, 0x2F, 0x57, 0x1C, 0x25,
	0x16, 0x1B, 0x0B, 0x18, 0x08, 0x0F, 0x59, 0x5D, 0x3F, 0x01, 0x38, 0x31,
	0x20, 0x11, 0x2B, 0x38, 0x54, 0x16, 0x1F, 0x35, 0x54, 0x0F, 0x14, 0x2F,
	0x08, 0x0A, 0x2B, 0x56, 0x1C, 0x3B, 0x20, 0x18, 0x08, 0x2A, 0x0D, 0x0E,
	0x31, 0x20, 0x53, 0x35, 0x00, 0x25, 0x14, 0x0D, 0x7A, 0x24, 0x0A, 0x5A,
	0x08, 0x20, 0x5A, 0x09, 0x06, 0x01, 0x38, 0x0A, 0x2C, 0x27, 0x08, 0x7A,
	0x5F, 0x19, 0x2C, 0x2F, 0x2C, 0x01, 0x4E, 0x01, 0x3F, 0x77, 0x59, 0x17,
	0x45, 0x2A, 0x24, 0x3E, 0x16, 0x3E, 0x09, 0x24, 0x55, 0x27, 0x38, 0x27,
	0x16, 0x39, 0x24, 0x41, 0x07, 0x11, 0x23, 0x0C, 0x34, 0x0A, 0x70, 0x06,
	0x10, 0x5E, 0x12, 0x32, 0x5F, 0x55, 0x01, 0x06, 0x0A, 0x04, 0x02, 0x1B,
	0x26, 0x04, 0x35, 0x04, 0x08, 0x2E, 0x2F, 0x5F, 0x58, 0x03, 0x03, 0x14,
	0x19, 0x34, 0x1C, 0x44, 0x76, 0x34, 0x07, 0x0D, 0x2E, 0x33, 0x5E, 0x58,
	0x1F, 0x28, 0x04, 0x26, 0x34, 0x58, 0x12, 0x2E, 0x26, 0x4A, 0x17, 0x3D,
	0x27, 0x16, 0x30, 0x23, 0x59, 0x20, 0x5F, 0x11, 0x16, 0x5B, 0x05, 0x3A,
	0x31, 0x24, 0x5B, 0x00, 0x0F, 0x57, 0x1F, 0x38, 0x08, 0x00, 0x22, 0x1A,
	0x25, 0x3A, 0x59, 0x34, 0x41, 0x11, 0x18, 0x55, 0x0D, 0x3E, 0x22, 0x37,
	0x5B, 0x09, 0x18, 0x39, 0x18, 0x55, 0x04, 0x26, 0x20, 0x2F, 0x21, 0x12,
	0x37, 0x02, 0x27, 0x5C, 0x19, 0x3B, 0x40, 0x2E, 0x2E, 0x11, 0x34, 0x24,
	0x0A, 0x1C, 0x39, 0x19, 0x05, 0x09, 0x21, 0x59, 0x0F, 0x0E, 0x73, 0x58,
	0x4E, 0x0B, 0x33, 0x18, 0x5A, 0x10, 0x1C, 0x3D, 0x38, 0x5C, 0x05, 0x1B,
	0x0E, 0x16, 0x3E, 0x16, 0x26, 0x3F, 0x15, 0x5D, 0x56, 0x21, 0x0A, 0x10,
	0x2A, 0x57, 0x5D, 0x2D, 0x3B, 0x1C, 0x10, 0x56, 0x44, 0x32, 0x54, 0x52,
	0x59, 0x05, 0x00, 0x3F, 0x52, 0x39, 0x29, 0x3A, 0x0F, 0x2F, 0x59, 0x04,
	0x07, 0x5E, 0x04, 0x01, 0x27, 0x11, 0x54, 0x13, 0x06, 0x08, 0x0B, 0x00,
	0x2A, 0x5B, 0x3D, 0x73, 0x18, 0x09, 0x41, 0x5F, 0x08, 0x47, 0x2B, 0x57,
	0x0C, 0x2F, 0x1E, 0x35, 0x1C, 0x2E, 0x32, 0x16, 0x31, 0x56, 0x18, 0x1A,
	0x5D, 0x2E, 0x0C, 0x19, 0x2F, 0x5C, 0x10, 0x3B, 0x44, 0x33, 0x00, 0x32,
	0x3A, 0x01, 0x2E, 0x15, 0x08, 0x58, 0x19, 0x0F, 0x1E, 0x27, 0x2F, 0x25,
	0x1A, 0x5B, 0x09, 0x2A, 0x1E, 0x16, 0x59, 0x35, 0x3B, 0x40, 0x1A, 0x19,
	0x50, 0x09, 0x2E, 0x16, 0x22, 0x56, 0x5C, 0x52, 0x33, 0x38, 0x16, 0x05,
	0x31, 0x72, 0x5E, 0x2E, 0x5B, 0x5F, 0x0A, 0x06, 0x10, 0x03, 0x44, 0x0D,
	0x5B, 0x09, 0x1A, 0x02, 0x1A, 0x5E, 0x0C, 0x00, 0x53, 0x2D, 0x29, 0x18,
	0x57, 0x58, 0x28, 0x59, 0x11, 0x09, 0x44, 0x09, 0x03, 0x50, 0x39, 0x26,
	0x04, 0x47, 0x56, 0x5C, 0x0D, 0x09, 0x3A, 0x57, 0x5B, 0x52, 0x33, 0x23,
	0x13, 0x0F, 0x0E, 0x15, 0x3E, 0x2A, 0x1A, 0x5B, 0x23, 0x5A, 0x09, 0x1B,
	0x3A, 0x72, 0x06, 0x52, 0x27, 0x0A, 0x15, 0x15, 0x36, 0x41, 0x03, 0x28,
	0x5D, 0x52, 0x2D, 0x13, 0x15, 0x55, 0x04, 0x19, 0x05, 0x03, 0x02, 0x0D,
	0x3E, 0x5D, 0x23, 0x5C, 0x00, 0x57, 0x01, 0x23, 0x1A, 0x0A, 0x18, 0x32,
	0x0D, 0x5A, 0x4A, 0x19, 0x38, 0x38, 0x05, 0x12, 0x56, 0x3D, 0x74, 0x34,
	0x59, 0x26, 0x1D, 0x33, 0x58, 0x2C, 0x59, 0x03, 0x1B, 0x19, 0x54, 0x23,
	0x32, 0x27, 0x0F, 0x16, 0x08, 0x0E, 0x16, 0x3B, 0x00, 0x5B, 0x58, 0x06,
	0x07, 0x37, 0x08, 0x3E, 0x00, 0x5F, 0x30, 0x21, 0x1F, 0x6D, 0x04, 0x02,
	0x14, 0x1E, 0x25, 0x39, 0x58, 0x05, 0x5F, 0x09, 0x3C, 0x52, 0x39, 0x40,
	0x17, 0x5D, 0x08, 0x1A, 0x0A, 0x0B, 0x2A, 0x13, 0x00, 0x5B, 0x77, 0x04,
	0x2E, 0x36, 0x44, 0x0E, 0x3F, 0x52, 0x1D, 0x07, 0x20, 0x23, 0x19, 0x16,
	0x1D, 0x01, 0x22, 0x02, 0x0C, 0x5D, 0x03, 0x09, 0x34, 0x29, 0x23, 0x17,
	0x29, 0x35, 0x5A, 0x5C, 0x10, 0x02, 0x2D, 0x1C, 0x58, 0x26, 0x05, 0x2E,
	0x56, 0x28, 0x21, 0x0E, 0x03, 0x18, 0x28, 0x37, 0x1A, 0x38, 0x01, 0x1C,
	0x12, 0x0A, 0x3B, 0x45, 0x53, 0x2E, 0x1F, 0x15, 0x03, 0x02, 0x09, 0x0F,
	0x15, 0x1A, 0x1E, 0x35, 0x0D, 0x26, 0x06, 0x52, 0x37, 0x2F, 0x2D, 0x1D,
	0x0E, 0x71, 0x0A, 0x3B, 0x25, 0x1F, 0x24, 0x3F, 0x1B, 0x08, 0x20, 0x35,
	0x18, 0x56, 0x1E, 0x3D, 0x21, 0x0F, 0x52, 0x58, 0x0D, 0x15, 0x1E, 0x18,
	0x0D, 0x24, 0x17, 0x03, 0x33, 0x59, 0x1B, 0x25, 0x5D, 0x2C, 0x21, 0x39,
	0x7A, 0x1E, 0x25, 0x3F, 0x5A, 0x04, 0x1F, 0x00, 0x0F, 0x19, 0x32, 0x07,
	0x27, 0x3C, 0x00, 0x37, 0x3A, 0x0B, 0x21, 0x1C, 0x24, 0x3C, 0x04, 0x21,
	0x33, 0x3B, 0x38, 0x39, 0x1C, 0x1F, 0x26, 0x09, 0x56, 0x23, 0x05, 0x12,
	0x5E, 0x0A, 0x3B, 0x11, 0x7B, 0x3F, 0x31, 0x2A, 0x11, 0x00, 0x23, 0x13,
	0x1C, 0x1A, 0x25, 0x18, 0x39, 0x41, 0x29, 0x31, 0x2D, 0x33, 0x02, 0x0E,
	0x12, 0x1C, 0x32, 0x06, 0x21, 0x01, 0x00, 0x14, 0x0B, 0x52, 0x00, 0x2B,
	0x22, 0x01, 0x05, 0x2F, 0x35, 0x33, 0x03, 0x3B, 0x2D, 0x1F, 0x31, 0x29,
	0x38, 0x1B, 0x35, 0x33, 0x5A, 0x09, 0x03, 0x01, 0x0B, 0x08, 0x3B, 0x0E,
	0x21, 0x12, 0x5E, 0x0F, 0x37, 0x20, 0x2E, 0x24, 0x08, 0x0A, 0x26, 0x27,
	0x1B, 0x0E, 0x34, 0x1C, 0x0C, 0x3A, 0x1F, 0x12, 0x1D, 0x17, 0x45, 0x2F,
	0x35, 0x1F, 0x39, 0x1A, 0x0E, 0x14, 0x34, 0x58, 0x03, 0x5F, 0x10, 0x28,
	0x04, 0x19, 0x5F, 0x29, 0x55, 0x13, 0x0C, 0x38, 0x34, 0x36, 0x00, 0x05,
	0x2F, 0x0C, 0x2B, 0x3B, 0x41, 0x59, 0x15, 0x00, 0x56, 0x3A, 0x3A, 0x17,
	0x5F, 0x10, 0x22, 0x1F, 0x74, 0x34, 0x50, 0x01, 0x33, 0x2D, 0x59, 0x1B,
	0x58, 0x31, 0x10, 0x24, 0x2A, 0x2D, 0x12, 0x70, 0x24, 0x22, 0x04, 0x3D,
	0x74, 0x16, 0x50, 0x16, 0x05, 0x21, 0x21, 0x4E, 0x3F, 0x5E, 0x07, 0x27,
	0x12, 0x00, 0x59, 0x24, 0x0E, 0x36, 0x22, 0x01, 0x37, 0x1E, 0x2F, 0x2C,
	0x3E, 0x3B, 0x5F, 0x1B, 0x05, 0x20, 0x2D, 0x3E, 0x17, 0x0B, 0x09, 0x1B,
	0x18, 0x50, 0x2B, 0x33, 0x2C, 0x0A, 0x14, 0x1D, 0x08, 0x15, 0x05, 0x24,
	0x5A, 0x32, 0x37, 0x20, 0x4E, 0x2F, 0x5F, 0x15, 0x54, 0x27, 0x0F, 0x1D,
	0x2F, 0x5B, 0x35, 0x06, 0x04, 0x13, 0x39, 0x28, 0x28, 0x1C, 0x69, 0x0A,
	0x12, 0x18, 0x2F, 0x3A, 0x23, 0x24, 0x5E, 0x3D, 0x28, 0x36, 0x20, 0x5B,
	0x26, 0x16, 0x1B, 0x30, 0x36, 0x1A, 0x37, 0x59, 0x52, 0x3E, 0x59, 0x37,
	0x3D, 0x59, 0x36, 0x26, 0x0D, 0x3B, 0x18, 0x0B, 0x52, 0x11, 0x39, 0x30,
	0x57, 0x0C, 0x6D, 0x29, 0x0D, 0x2D, 0x53, 0x7A, 0x1E, 0x2D, 0x1C, 0x13,
	0x18, 0x3F, 0x39, 0x00, 0x03, 0x3B, 0x07, 0x28, 0x29, 0x53, 0x14, 0x05,
	0x0B, 0x29, 0x26, 0x7B, 0x34, 0x50, 0x16, 0x1C, 0x14, 0x1C, 0x54, 0x58,
	0x27, 0x03, 0x39, 0x28, 0x5F, 0x19, 0x07, 0x54, 0x56, 0x16, 0x5C, 0x20,
	0x5B, 0x08, 0x0D, 0x26, 0x7B, 0x16, 0x12, 0x5D, 0x32, 0x27, 0x26, 0x11,
	0x26, 0x2E, 0x36, 0x0E, 0x18, 0x1E, 0x2A, 0x05, 0x16, 0x54, 0x5B, 0x52,
	0x2C, 0x28, 0x11, 0x17, 0x59, 0x00, 0x3E, 0x07, 0x37, 0x13, 0x3B, 0x0E,
	0x52, 0x06, 0x5D, 0x26, 0x47, 0x26, 0x04, 0x04, 0x38, 0x05, 0x24, 0x14,
	0x40, 0x70, 0x06, 0x51, 0x07, 0x1B, 0x2B, 0x2D, 0x27, 0x41, 0x08, 0x6D,
	0x47, 0x04, 0x1F, 0x04, 0x11, 0x08, 0x56, 0x3D, 0x11, 0x73, 0x1F, 0x53,
	0x14, 0x2C, 0x2E, 0x47, 0x02, 0x3C, 0x28, 0x34, 0x1A, 0x31, 0x00, 0x5E,
	0x37, 0x1D, 0x29, 0x1B, 0x20, 0x0E, 0x3C, 0x0D, 0x3F, 0x08, 0x7B, 0x06,
	0x39, 0x1B, 0x58, 0x10, 0x1B, 0x1B, 0x41, 0x24, 0x6D, 0x1D, 0x0B, 0x39,
	0x5D, 0x72, 0x0E, 0x07, 0x14, 0x0F, 0x2B, 0x55, 0x09, 0x5F, 0x06, 0x06,
	0x47, 0x0A, 0x0C, 0x01, 0x27, 0x5F, 0x07, 0x0F, 0x38, 0x69, 0x04, 0x23,
	0x14, 0x40, 0x33, 0x14, 0x57, 0x14, 0x2D, 0x00, 0x07, 0x4E, 0x59, 0x0A,
	0x28, 0x00, 0x05, 0x01, 0x12, 0x23, 0x25, 0x31, 0x2C, 0x26, 0x69, 0x08,
	0x52, 0x18, 0x12, 0x29, 0x54, 0x04, 0x41, 0x11, 0x03, 0x36, 0x13, 0x5A,
	0x1D, 0x33, 0x1F, 0x0F, 0x23, 0x44, 0x34, 0x5D, 0x02, 0x57, 0x11, 0x13,
	0x18, 0x2B, 0x27, 0x5A, 0x0E, 0x0F, 0x59, 0x5A, 0x29, 0x04, 0x55, 0x05,
	0x56, 0x19, 0x2D, 0x5E, 0x17, 0x3B, 0x3D, 0x70, 0x3F, 0x04, 0x08, 0x18,
	0x2F, 0x02, 0x36, 0x22, 0x3D, 0x74, 0x43, 0x25, 0x41, 0x0D, 0x13, 0x43,
	0x58, 0x36, 0x05, 0x7A, 0x0E, 0x14, 0x01, 0x22, 0x7A, 0x3E, 0x53, 0x25,
	0x03, 0x11, 0x01, 0x27, 0x07, 0x1F, 0x69, 0x25, 0x05, 0x18, 0x03, 0x30,
	0x5B, 0x2E, 0x18, 0x5F, 0x37, 0x39, 0x2E, 0x1B, 0x40, 0x27, 0x55, 0x57,
	0x5B, 0x03, 0x27, 0x2D, 0x08, 0x5F, 0x52, 0x77, 0x2E, 0x03, 0x57, 0x19,
	0x21, 0x3E, 0x39, 0x05, 0x3E, 0x00, 0x18, 0x2F, 0x26, 0x1F, 0x77, 0x35,
	0x06, 0x03, 0x44, 0x24, 0x34, 0x2D, 0x2B, 0x59, 0x74, 0x15, 0x0D, 0x38,
	0x52, 0x7A, 0x0D, 0x2C, 0x3B, 0x08, 0x72, 0x55, 0x2D, 0x18, 0x5C, 0x07,
	0x20, 0x50, 0x00, 0x2C, 0x2E, 0x1C, 0x56, 0x0A, 0x39, 0x18, 0x02, 0x15,
	0x59, 0x59, 0x16, 0x20, 0x22, 0x02, 0x05, 0x36, 0x04, 0x07, 0x41, 0x00,
	0x7A, 0x16, 0x00, 0x25, 0x07, 0x32, 0x0A, 0x14, 0x07, 0x26, 0x09, 0x24,
	0x31, 0x36, 0x11, 0x07, 0x1D, 0x2C, 0x2C, 0x3B, 0x2A, 0x2A, 0x56, 0x3D,
	0x26, 0x23, 0x06, 0x04, 0x5C, 0x23, 0x0C, 0x5B, 0x15, 0x36, 0x19, 0x0F,
	0x5E, 0x27, 0x18, 0x1D, 0x7A, 0x29, 0x00, 0x57, 0x2E, 0x11, 0x5F, 0x03,
	0x02, 0x52, 0x23, 0x47, 0x50, 0x04, 0x29, 0x08, 0x15, 0x37, 0x05, 0x5D,
	0x72, 0x2E, 0x34, 0x08, 0x5A, 0x14, 0x06, 0x19, 0x1E, 0x27, 0x07, 0x03,
	0x07, 0x5F, 0x1D, 0x35, 0x2B, 0x15, 0x05, 0x28, 0x30, 0x5B, 0x04, 0x02,
	0x40, 0x03, 0x21, 0x2B, 0x08, 0x40, 0x15, 0x0F, 0x23, 0x14, 0x59, 0x0C,
	0x47, 0x12, 0x5C, 0x3E, 0x37, 0x35, 0x34, 0x23, 0x0D, 0x1B, 0x59, 0x0F,
	0x22, 0x20, 0x2E, 0x55, 0x50, 0x22, 0x3B, 0x14, 0x36, 0x10, 0x08, 0x1C,
	0x35, 0x26, 0x0E, 0x00, 0x0E, 0x69, 0x5B, 0x00, 0x5A, 0x0C, 0x05, 0x2A,
	0x56, 0x00, 0x0D, 0x37, 0x0E, 0x54, 0x14, 0x08, 0x0C, 0x2B, 0x4E, 0x0A,
	0x11, 0x06, 0x5A, 0x13, 0x29, 0x1A, 0x20, 0x0B, 0x32, 0x45, 0x5C, 0x14,
	0x04, 0x0A, 0x39, 0x2D, 0x0E, 0x0B, 0x17, 0x5B, 0x27, 0x0C, 0x5A, 0x00,
	0x5B, 0x2D, 0x7B, 0x5B, 0x23, 0x5D, 0x44, 0x13, 0x39, 0x09, 0x2D, 0x40,
	0x74, 0x26, 0x13, 0x34, 0x24, 0x6D, 0x0A, 0x31, 0x3F, 0x38, 0x26, 0x02,
	0x29, 0x59, 0x0D, 0x07, 0x03, 0x59, 0x5D, 0x5C, 0x20, 0x3C, 0x54, 0x5C,
	0x27, 0x28, 0x3B, 0x13, 0x3A, 0x05, 0x03, 0x1A, 0x00, 0x5C, 0x08, 0x30,
	0x24, 0x59, 0x45, 0x5B, 0x24, 0x04, 0x2A, 0x39, 0x0D, 0x75, 0x04, 0x57,
	0x5F, 0x1F, 0x0A, 0x27, 0x08, 0x2F, 0x1F, 0x0E, 0x22, 0x50, 0x5D, 0x2D,
	0x29, 0x5F, 0x57, 0x3B, 0x25, 0x70, 0x16, 0x39, 0x14, 0x5A, 0x7A, 0x07,
	0x58, 0x22, 0x03, 0x10, 0x0D, 0x27, 0x0C, 0x33, 0x06, 0x15, 0x4A, 0x37,
	0x32, 0x2E, 0x54, 0x03, 0x26, 0x33, 0x12, 0x1E, 0x10, 0x28, 0x5E, 0x13,
	0x5C, 0x31, 0x06, 0x29, 0x0A, 0x04, 0x31, 0x16, 0x08, 0x1A, 0x08, 0x4A,
	0x5B, 0x0C, 0x70, 0x5D, 0x2D, 0x1C, 0x0E, 0x09, 0x34, 0x13, 0x26, 0x28,
	0x23, 0x3B, 0x4E, 0x0A, 0x3C, 0x16, 0x14, 0x4E, 0x17, 0x40, 0x32, 0x20,
	0x16, 0x5A, 0x0A, 0x71, 0x5F, 0x35, 0x0C, 0x12, 0x27, 0x34, 0x32, 0x0F,
	0x40, 0x75, 0x21, 0x39, 0x18, 0x02, 0x10, 0x54, 0x19, 0x1D, 0x06, 0x10,
	0x03, 0x52, 0x22, 0x28, 0x3A, 0x1F, 0x51, 0x14, 0x06, 0x1A, 0x38, 0x19,
	0x21, 0x29, 0x34, 0x5F, 0x07, 0x2A, 0x2C, 0x0B, 0x5E, 0x4E, 0x08, 0x29,
	0x03, 0x1A, 0x2F, 0x57, 0x05, 0x69, 0x27, 0x50, 0x08, 0x1C, 0x76, 0x59,
	0x08, 0x1D, 0x52, 0x76, 0x5E, 0x54, 0x3A, 0x08, 0x0F, 0x3C, 0x27, 0x0B,
	0x52, 0x0C, 0x15, 0x17, 0x5A, 0x12, 0x3B, 0x20, 0x19, 0x06, 0x05, 0x2B,
	0x3B, 0x55, 0x0C, 0x38, 0x70, 0x01, 0x04, 0x3B, 0x27, 0x10, 0x06, 0x57,
	0x5A, 0x3A, 0x36, 0x43, 0x52, 0x5D, 0x03, 0x69, 0x20, 0x2F, 0x59, 0x1C,
	0x18, 0x0A, 0x55, 0x24, 0x0A, 0x17, 0x1E, 0x37, 0x02, 0x11, 0x21, 0x24,
	0x00, 0x39, 0x0A, 0x24, 0x1E, 0x14, 0x14, 0x2C, 0x2C, 0x55, 0x18, 0x34,
	0x00, 0x28, 0x3C, 0x00, 0x45, 0x44, 0x33, 0x5F, 0x06, 0x57, 0x0D, 0x11,
	0x24, 0x36, 0x23, 0x0D, 0x23, 0x09, 0x2C, 0x1C, 0x19, 0x6D, 0x3B, 0x57,
	0x19, 0x0F, 0x05, 0x08, 0x0D, 0x3A, 0x53, 0x25, 0x1B, 0x2D, 0x57, 0x5F,
	0x26, 0x47, 0x19, 0x01, 0x05, 0x06, 0x27, 0x0B, 0x36, 0x52, 0x00, 0x39,
	0x16, 0x5B, 0x08, 0x3A, 0x23, 0x53, 0x25, 0x02, 0x07, 0x02, 0x13, 0x18,
	0x59, 0x1B, 0x04, 0x39, 0x08, 0x11, 0x2A, 0x3D, 0x07, 0x1E, 0x33, 0x73,
	0x43, 0x15, 0x2D, 0x07, 0x23, 0x23, 0x02, 0x45, 0x0E, 0x2A, 0x3B, 0x10,
	0x45, 0x2F, 0x74, 0x5B, 0x4E, 0x1E, 0x26, 0x2D, 0x16, 0x03, 0x18, 0x40,
	0x09, 0x18, 0x13, 0x06, 0x06, 0x75, 0x3E, 0x0E, 0x3B, 0x03, 0x06, 0x47,
	0x59, 0x3E, 0x01, 0x07, 0x35, 0x2E, 0x39, 0x07, 0x26, 0x58, 0x2B, 0x36,
	0x13, 0x3A, 0x0B, 0x02, 0x41, 0x44, 0x20, 0x5F, 0x22, 0x02, 0x11, 0x38,
	0x39, 0x2E, 0x27, 0x0E, 0x32, 0x38, 0x37, 0x0C, 0x58, 0x36, 0x0E, 0x51,
	0x03, 0x23, 0x12, 0x1B, 0x04, 0x2F, 0x20, 0x0D, 0x3A, 0x18, 0x3C, 0x25,
	0x2B, 0x38, 0x15, 0x14, 0x1D, 0x2F, 0x2B, 0x29, 0x01, 0x26, 0x69, 0x0E,
	0x19, 0x58, 0x5A, 0x14, 0x3C, 0x17, 0x07, 0x00, 0x76, 0x0F, 0x12, 0x0A,
	0x03, 0x1A, 0x01, 0x10, 0x3D, 0x12, 0x37, 0x0A, 0x03, 0x22, 0x18, 0x75,
	0x0F, 0x2F, 0x2C, 0x53, 0x34, 0x23, 0x2B, 0x3D, 0x18, 0x24, 0x09, 0x59,
	0x0F, 0x3B, 0x15, 0x38, 0x16, 0x1E, 0x3C, 0x0E, 0x59, 0x13, 0x41, 0x0F,
	0x7A, 0x14, 0x0D, 0x5D, 0x06, 0x3A, 0x1C, 0x36, 0x5F, 0x5D, 0x34, 0x14,
	0x52, 0x21, 0x0E, 0x74, 0x0D, 0x00, 0x18, 0x2C, 0x0E, 0x0E, 0x03, 0x16,
	0x1C, 0x04, 0x34, 0x39, 0x24, 0x2E, 0x7B, 0x09, 0x2F, 0x17, 0x19, 0x1A,
	0x0D, 0x05, 0x04, 0x01, 0x72, 0x1A, 0x07, 0x2A, 0x01, 0x31, 0x5B, 0x22,
	0x58, 0x53, 0x75, 0x43, 0x03, 0x2C, 0x20, 0x20, 0x20, 0x12, 0x27, 0x1D,
	0x7B, 0x04, 0x13, 0x5A, 0x5E, 0x33, 0x20, 0x51, 0x24, 0x0E, 0x74, 0x59,
	0x02, 0x18, 0x3C, 0x25, 0x24, 0x0E, 0x5A, 0x44, 0x34, 0x39, 0x4E, 0x39,
	0x5E, 0x7B, 0x58, 0x12, 0x1B, 0x1E, 0x23, 0x2D, 0x12, 0x41, 0x13, 0x2F,
	0x5B, 0x2D, 0x5E, 0x5C, 0x26, 0x0A, 0x08, 0x5F, 0x0D, 0x7A, 0x5B, 0x04,
	0x00, 0x3B, 0x70, 0x0B, 0x03, 0x2D, 0x1B, 0x0D, 0x1A, 0x4E, 0x28, 0x02,
	0x14, 0x0F, 0x2C, 0x0F, 0x28, 0x21, 0x3C, 0x2A, 0x3C, 0x3C, 0x0B, 0x08,
	0x0F, 0x08, 0x04, 0x13, 0x34, 0x4E, 0x06, 0x5B, 0x38, 0x43, 0x0E, 0x00,
	0x0D, 0x30, 0x01, 0x39, 0x0C, 0x1E, 0x0D, 0x59, 0x58, 0x16, 0x0A, 0x36,
	0x24, 0x38, 0x27, 0x0D, 0x74, 0x38, 0x15, 0x0B, 0x08, 0x31, 0x54, 0x16,
	0x17, 0x02, 0x37, 0x1F, 0x3B, 0x03, 0x23, 0x07, 0x1F, 0x37, 0x05, 0x5E,
	0x69, 0x2F, 0x22, 0x21, 0x5B, 0x3B, 0x5A, 0x25, 0x1D, 0x38, 0x69, 0x28,
	0x0F, 0x59, 0x5C, 0x12, 0x18, 0x52, 0x19, 0x5E, 0x69, 0x2D, 0x03, 0x1B,
	0x0F, 0x33, 0x1D, 0x3B, 0x16, 0x08, 0x30, 0x0E, 0x15, 0x45, 0x0E, 0x09,
	0x27, 0x18, 0x1B, 0x59, 0x1B, 0x0E, 0x0A, 0x5B, 0x19, 0x34, 0x20, 0x26,
	0x21, 0x28, 0x05, 0x47, 0x19, 0x56, 0x24, 0x76, 0x2B, 0x12, 0x0F, 0x0A,
	0x0C, 0x16, 0x2E, 0x1F, 0x18, 0x6D, 0x2F, 0x57, 0x19, 0x3C, 0x18, 0x19,
	0x39, 0x45, 0x5C, 0x70, 0x47, 0x2E, 0x04, 0x3A, 0x21, 0x47, 0x3B, 0x5C,
	0x1A, 0x24, 0x5C, 0x27, 0x41, 0x26, 0x10, 0x07, 0x06, 0x5B, 0x27, 0x08,
	0x3D, 0x33, 0x38, 0x25, 0x17, 0x5B, 0x0D, 0x21, 0x2C, 0x24, 0x0D, 0x0F,
	0x45, 0x1E, 0x09, 0x36, 0x12, 0x3B, 0x5B, 0x06, 0x0E, 0x15, 0x41, 0x0F,
	0x27, 0x54, 0x37, 0x1D, 0x25, 0x2C, 0x5B, 0x4A, 0x1E, 0x1C, 0x72, 0x24,
	0x13, 0x45, 0x3D, 0x26, 0x15, 0x03, 0x19, 0x0A, 0x12, 0x1D, 0x27, 0x03,
	0x53, 0x74, 0x18, 0x11, 0x1C, 0x02, 0x21, 0x01, 0x0F, 0x56, 0x3F, 0x34,
	0x39, 0x07, 0x29, 0x44, 0x33, 0x06, 0x58, 0x23, 0x1D, 0x2B, 0x5D, 0x50,
	0x5D, 0x24, 0x36, 0x5B, 0x32, 0x25, 0x18, 0x2C, 0x24, 0x09, 0x03, 0x22,
	0x23, 0x47, 0x4E, 0x0C, 0x08, 0x77, 0x1A, 0x53, 0x1E, 0x23, 0x28, 0x54,
	0x58, 0x3D, 0x0F, 0x1A, 0x58, 0x52, 0x2D, 0x19, 0x18, 0x38, 0x57, 0x38,
	0x2F, 0x6D, 0x1E, 0x34, 0x36, 0x40, 0x6D, 0x55, 0x18, 0x25, 0x05, 0x37,
	0x24, 0x14, 0x3B, 0x2A, 0x24, 0x07, 0x33, 0x03, 0x59, 0x17, 0x18, 0x35,
	0x3E, 0x11, 0x04, 0x59, 0x13, 0x5F, 0x0A, 0x6D, 0x02, 0x4A, 0x00, 0x3F,
	0x26, 0x0A, 0x24, 0x1A, 0x22, 0x6D, 0x35, 0x52, 0x02, 0x12, 0x69, 0x09,
	0x07, 0x21, 0x21, 0x69, 0x0D, 0x29, 0x1F, 0x29, 0x7A, 0x03, 0x3B, 0x27,
	0x0D, 0x06, 0x5A, 0x15, 0x0B, 0x32, 0x38, 0x55, 0x59, 0x20, 0x1F, 0x06,
	0x0E, 0x53, 0x5A, 0x04, 0x15, 0x34, 0x29, 0x1B, 0x5B, 0x2E, 0x0E, 0x59,
	0x03, 0x3B, 0x33, 0x0F, 0x36, 0x58, 0x1D, 0x12, 0x1D, 0x30, 0x59, 0x05,
	0x00, 0x28, 0x09, 0x23, 0x2C, 0x70, 0x09, 0x0C, 0x09, 0x3A, 0x6D, 0x3B,
	0x55, 0x1E, 0x3C, 0x30, 0x24, 0x27, 0x0F, 0x33, 0x36, 0x22, 0x59, 0x1F,
	0x32, 0x28, 0x18, 0x12, 0x34, 0x1E, 0x04, 0x23, 0x37, 0x17, 0x44, 0x23,
	0x5D, 0x3B, 0x02, 0x0D, 0x36, 0x01, 0x55, 0x18, 0x0D, 0x6D, 0x2F, 0x50,
	0x18, 0x33, 0x76, 0x22, 0x39, 0x02, 0x13, 0x26, 0x36, 0x31, 0x1E, 0x11,
	0x7A, 0x36, 0x11, 0x59, 0x21, 0x76, 0x5E, 0x29, 0x16, 0x20, 0x73, 0x59,
	0x35, 0x23, 0x2E, 0x24, 0x38, 0x35, 0x24, 0x25, 0x0D, 0x3A, 0x54, 0x3F,
	0x1E, 0x69, 0x28, 0x50, 0x2F, 0x59, 0x24, 0x24, 0x16, 0x22, 0x1D, 0x69,
	0x09, 0x2A, 0x14, 0x24, 0x32, 0x1D, 0x0C, 0x1A, 0x5F, 0x76, 0x5A, 0x55,
	0x0C, 0x32, 0x37, 0x01, 0x38, 0x2D, 0x09, 0x74, 0x05, 0x4E, 0x2B, 0x58,
	0x7A, 0x47, 0x03, 0x29, 0x3B, 0x7B, 0x43, 0x52, 0x5A, 0x05, 0x38, 0x07,
	0x34, 0x29, 0x33, 0x34, 0x22, 0x38, 0x1B, 0x44, 0x76, 0x54, 0x56, 0x26,
	0x01, 0x2C, 0x15, 0x4E, 0x0B, 0x01, 0x1A, 0x1F, 0x19, 0x5A, 0x2E, 0x14,
	0x3F, 0x13, 0x23, 0x2C, 0x27, 0x24, 0x0F, 0x07, 0x07, 0x0F, 0x2A, 0x03,
	0x18, 0x1B, 0x70, 0x04, 0x02, 0x27, 0x0A, 0x36, 0x55, 0x57, 0x38, 0x26,
	0x71, 0x2A, 0x24, 0x45, 0x29, 0x3B, 0x55, 0x50, 0x2D, 0x1D, 0x7B, 0x5A,
	0x16, 0x20, 0x44, 0x30, 0x58, 0x0A, 0x07, 0x2F, 0x72, 0x18, 0x2A, 0x0B,
	0x0E, 0x7B, 0x43, 0x06, 0x2A, 0x3A, 0x2C, 0x34, 0x04, 0x59, 0x52, 0x75,
	0x01, 0x39, 0x24, 0x38, 0x18, 0x5C, 0x56, 0x2A, 0x1D, 0x2E, 0x5D, 0x39,
	0x00, 0x23, 0x04, 0x3A, 0x58, 0x59, 0x19, 0x07, 0x02, 0x33, 0x1D, 0x13,
	0x30, 0x1E, 0x56, 0x1A, 0x11, 0x12, 0x05, 0x19, 0x18, 0x02, 0x14, 0x58,
	0x34, 0x21, 0x2F, 0x29, 0x35, 0x59, 0x34, 0x33, 0x2B, 0x55, 0x37, 0x18,
	0x0D, 0x17, 0x1A, 0x56, 0x56, 0x07, 0x20, 0x43, 0x2A, 0x38, 0x5D, 0x27,
	0x23, 0x37, 0x3A, 0x2E, 0x2F, 0x43, 0x00, 0x39, 0x08, 0x71, 0x5B, 0x0D,
	0x1B, 0x1E, 0x15, 0x22, 0x24, 0x06, 0x1F, 0x7A, 0x5B, 0x59, 0x14, 0x08,
	0x7A, 0x29, 0x17, 0x1C, 0x26, 0x2F, 0x3A, 0x07, 0x25, 0x28, 0x0C, 0x55,
	0x2D, 0x1A, 0x1F, 0x0F, 0x14, 0x0D, 0x0B, 0x07, 0x05, 0x1B, 0x52, 0x17,
	0x1E, 0x2A, 0x0B, 0x0E, 0x45, 0x5A, 0x11, 0x5A, 0x02, 0x18, 0x3F, 0x17,
	0x03, 0x51, 0x5C, 0x5F, 0x17, 0x01, 0x2B, 0x39, 0x3E, 0x7A, 0x1D, 0x25,
	0x21, 0x0A, 0x26, 0x21, 0x13, 0x1B, 0x26, 0x0E, 0x59, 0x06, 0x01, 0x23,
	0x76, 0x3F, 0x37, 0x26, 0x31, 0x73, 0x3A, 0x06, 0x3E, 0x09, 0x08, 0x18,
	0x0C, 0x19, 0x25, 0x30, 0x0F, 0x17, 0x0B, 0x3B, 0x2C, 0x03, 0x30, 0x3E,
	0x0A, 0x00, 0x01, 0x59, 0x1C, 0x5C, 0x25, 0x5F, 0x00, 0x5F, 0x01, 0x16,
	0x5B, 0x39, 0x5F, 0x39, 0x7B, 0x29, 0x50, 0x41, 0x5F, 0x76, 0x09, 0x14,
	0x04, 0x0E, 0x1A, 0x36, 0x1B, 0x0F, 0x25, 0x18, 0x28, 0x2A, 0x1F, 0x09,
	0x74, 0x5F, 0x19, 0x04, 0x21, 0x2A, 0x5C, 0x07, 0x23, 0x26, 0x0C, 0x09,
	0x34, 0x07, 0x28, 0x09, 0x09, 0x26, 0x5F, 0x58, 0x7B, 0x25, 0x31, 0x18,
	0x03, 0x23, 0x5D, 0x11, 0x45, 0x22, 0x76, 0x34, 0x31, 0x5D, 0x0D, 0x27,
	0x28, 0x3B, 0x0A, 0x0A, 0x2C, 0x08, 0x08, 0x17, 0x31, 0x7A, 0x2B, 0x16,
	0x29, 0x11, 0x1A, 0x58, 0x54, 0x3A, 0x5B, 0x2C, 0x3B, 0x33, 0x0D, 0x08,
	0x75, 0x38, 0x50, 0x17, 0x5B, 0x29, 0x23, 0x26, 0x0C, 0x11, 0x3A, 0x1E,
	0x06, 0x1D, 0x1D, 0x2B, 0x34, 0x10, 0x56, 0x5E, 0x14, 0x02, 0x18, 0x07,
	0x5C, 0x28, 0x03, 0x0D, 0x3B, 0x33, 0x0E, 0x2A, 0x2E, 0x3F, 0x23, 0x71,
	0x47, 0x15, 0x09, 0x12, 0x7A, 0x5E, 0x39, 0x14, 0x1A, 0x74, 0x22, 0x50,
	0x1E, 0x39, 0x76, 0x5E, 0x17, 0x00, 0x5E, 0x14, 0x47, 0x26, 0x0F, 0x58,
	0x7B, 0x1B, 0x17, 0x00, 0x0A, 0x7B, 0x5C, 0x30, 0x41, 0x1B, 0x38, 0x43,
	0x2F, 0x2B, 0x5E, 0x7B, 0x1F, 0x20, 0x28, 0x40, 0x75, 0x0E, 0x18, 0x20,
	0x13, 0x70, 0x2B, 0x00, 0x0B, 0x18, 0x12, 0x14, 0x16, 0x5D, 0x5B, 0x12,
	0x3F, 0x25, 0x59, 0x2C, 0x76, 0x2B, 0x37, 0x5B, 0x39, 0x7B, 0x39, 0x53,
	0x3C, 0x00, 0x2A, 0x39, 0x05, 0x02, 0x03, 0x1B, 0x1E, 0x2F, 0x18, 0x5A,
	0x20, 0x05, 0x02, 0x0B, 0x22, 0x10, 0x2A, 0x00, 0x2C, 0x29, 0x30, 0x5E,
	0x2D, 0x24, 0x3C, 0x76, 0x24, 0x0B, 0x0C, 0x33, 0x12, 0x1D, 0x18, 0x28,
	0x3C, 0x69, 0x5A, 0x57, 0x57, 0x05, 0x30, 0x21, 0x56, 0x3A, 0x5F, 0x21,
	0x20, 0x17, 0x38, 0x31, 0x14, 0x1A, 0x52, 0x3A, 0x3E, 0x0A, 0x15, 0x07,
	0x17, 0x32, 0x38, 0x2E, 0x14, 0x5C, 0x05, 0x08, 0x5B, 0x33, 0x0D, 0x28,
	0x08, 0x03, 0x08, 0x38, 0x23, 0x70, 0x16, 0x20, 0x0F, 0x0D, 0x17, 0x20,
	0x2B, 0x18, 0x53, 0x36, 0x0E, 0x17, 0x08, 0x12, 0x27, 0x02, 0x39, 0x00,
	0x31, 0x31, 0x5D, 0x24, 0x28, 0x0F, 0x38, 0x0B, 0x13, 0x20, 0x1F, 0x36,
	0x5B, 0x57, 0x2B, 0x05, 0x30, 0x1B, 0x33, 0x18, 0x23, 0x2B, 0x5C, 0x33,
	0x3B, 0x21, 0x2F, 0x58, 0x59, 0x0F, 0x08, 0x18, 0x18, 0x2F, 0x29, 0x23,
	0x31, 0x5F, 0x1B, 0x59, 0x5D, 0x13, 0x5F, 0x0A, 0x5F, 0x1A, 0x31, 0x1F,
	0x19, 0x5C, 0x5A, 0x28, 0x28, 0x53, 0x17, 0x0F, 0x12, 0x5B, 0x4E, 0x5E,
	0x1C, 0x2D, 0x2B, 0x2D, 0x1A, 0x44, 0x3A, 0x55, 0x4E, 0x3A, 0x2D, 0x7A,
	0x21, 0x10, 0x57, 0x0D, 0x32, 0x23, 0x17, 0x06, 0x31, 0x7B, 0x43, 0x3B,
	0x24, 0x5C, 0x13, 0x0E, 0x16, 0x58, 0x24, 0x7A, 0x54, 0x05, 0x06, 0x27,
	0x14, 0x00, 0x3B, 0x3B, 0x02, 0x76, 0x09, 0x35, 0x04, 0x1C, 0x74, 0x08,
	0x2B, 0x57, 0x00, 0x7A, 0x1F, 0x33, 0x25, 0x58, 0x7B, 0x3E, 0x28, 0x25,
	0x2A, 0x2E, 0x58, 0x17, 0x20, 0x06, 0x2C, 0x26, 0x27, 0x36, 0x2D, 0x0A,
	0x00, 0x52, 0x5D, 0x2E, 0x75, 0x5E, 0x4A, 0x17, 0x3D, 0x0A, 0x1F, 0x37,
	0x5C, 0x09, 0x75, 0x5B, 0x52, 0x3B, 0x3F, 0x73, 0x36, 0x4A, 0x26, 0x33,
	0x71, 0x0A, 0x23, 0x28, 0x52, 0x13, 0x58, 0x00, 0x09, 0x5A, 0x75, 0x47,
	0x56, 0x22, 0x58, 0x30, 0x5F, 0x2A, 0x04, 0x3D, 0x25, 0x55, 0x33, 0x03,
	0x5F, 0x29, 0x08, 0x2D, 0x3A, 0x5A, 0x71, 0x09, 0x0A, 0x41, 0x13, 0x38,
	0x1A, 0x02, 0x00, 0x03, 0x00, 0x5E, 0x39, 0x5C, 0x2D, 0x74, 0x34, 0x55,
	0x16, 0x58, 0x73, 0x0A, 0x11, 0x1C, 0x5D, 0x27, 0x54, 0x28, 0x2D, 0x0A,
	0x75, 0x0E, 0x25, 0x57, 0x1C, 0x76, 0x3D, 0x08, 0x0B, 0x58, 0x38, 0x1A,
	0x0C, 0x05, 0x52, 0x2F, 0x5E, 0x1B, 0x5B, 0x23, 0x33, 0x3B, 0x13, 0x24,
	0x2D, 0x37, 0x5F, 0x54, 0x08, 0x27, 0x7A, 0x3D, 0x39, 0x58, 0x58, 0x74,
	0x35, 0x39, 0x21, 0x00, 0x21, 0x25, 0x0B, 0x58, 0x5A, 0x23, 0x26, 0x0B,
	0x0D, 0x08, 0x09, 0x03, 0x4A, 0x41, 0x02, 0x18, 0x1C, 0x50, 0x45, 0x00,
	0x00, 0x15, 0x18, 0x3E, 0x08, 0x1A, 0x14, 0x12, 0x3E, 0x13, 0x73, 0x26,
	0x08, 0x16, 0x1A, 0x0F, 0x0A, 0x56, 0x04, 0x1D, 0x12, 0x23, 0x25, 0x16,
	0x0E, 0x74, 0x18, 0x35, 0x0B, 0x07, 0x12, 0x58, 0x51, 0x1E, 0x1A, 0x1A,
	0x3D, 0x0B, 0x19, 0x5C, 0x2B, 0x1E, 0x2B, 0x04, 0x24, 0x27, 0x47, 0x0B,
	0x3A, 0x0A, 0x12, 0x26, 0x52, 0x3E, 0x3E, 0x01, 0x05, 0x16, 0x37, 0x53,
	0x3A, 0x3B, 0x0B, 0x58, 0x52, 0x36, 0x3C, 0x0F, 0x16, 0x1F, 0x3B, 0x5F,
	0x18, 0x28, 0x5C, 0x05, 0x3F, 0x28, 0x1D, 0x31, 0x25, 0x26, 0x58, 0x0B,
	0x05, 0x36, 0x04, 0x0E, 0x57, 0x59, 0x14, 0x34, 0x11, 0x21, 0x5A, 0x2E,
	0x3B, 0x03, 0x3D, 0x1D, 0x26, 0x3F, 0x00, 0x0B, 0x5C, 0x24, 0x22, 0x05,
	0x56, 0x40, 0x27, 0x2E, 0x2E, 0x5F, 0x09, 0x06, 0x38, 0x11, 0x5F, 0x5D,
	0x0C, 0x08, 0x4A, 0x1A, 0x2D, 0x2C, 0x47, 0x14, 0x38, 0x01, 0x28, 0x25,
	0x05, 0x25, 0x44, 0x2E, 0x18, 0x58, 0x24, 0x09, 0x1A, 0x5A, 0x57, 0x3E,
	0x20, 0x69, 0x01, 0x25, 0x03, 0x5F, 0x70, 0x27, 0x53, 0x56, 0x1E, 0x77,
	0x1A, 0x59, 0x56, 0x1F, 0x77, 0x09, 0x58, 0x3E, 0x0F, 0x13, 0x59, 0x4E,
	0x24, 0x0E, 0x07, 0x1A, 0x19, 0x1B, 0x44, 0x34, 0x09, 0x53, 0x1C, 0x03,
	0x35, 0x43, 0x2E, 0x00, 0x1D, 0x00, 0x5E, 0x0F, 0x04, 0x28, 0x25, 0x43,
	0x0B, 0x1B, 0x44, 0x32, 0x3A, 0x02, 0x00, 0x44, 0x21, 0x02, 0x1B, 0x3B,
	0x1D, 0x14, 0x1B, 0x50, 0x0C, 0x2C, 0x26, 0x0B, 0x0A, 0x16, 0x2E, 0x27,
	0x5D, 0x59, 0x56, 0x1B, 0x73, 0x24, 0x0F, 0x26, 0x03, 0x0D, 0x19, 0x2D,
	0x20, 0x27, 0x3B, 0x34, 0x19, 0x01, 0x0A, 0x0F, 0x1B, 0x16, 0x57, 0x32,
	0x76, 0x3E, 0x15, 0x56, 0x32, 0x73, 0x15, 0x38, 0x19, 0x5C, 0x16, 0x28,
	0x53, 0x1A, 0x44, 0x72, 0x5E, 0x55, 0x08, 0x19, 0x0A, 0x01, 0x52, 0x0B,
	0x20, 0x12, 0x5B, 0x02, 0x3A, 0x5E, 0x37, 0x04, 0x58, 0x1C, 0x5C, 0x26,
	0x23, 0x38, 0x1F, 0x2C, 0x0E, 0x59, 0x32, 0x21, 0x04, 0x13, 0x5C, 0x37,
	0x3A, 0x0C, 0x3B, 0x20, 0x0F, 0x1C, 0x59, 0x30, 0x1D, 0x26, 0x3C, 0x1C,
	0x00, 0x24, 0x57, 0x05, 0x1D, 0x74, 0x5E, 0x23, 0x1F, 0x5A, 0x75, 0x36,
	0x51, 0x57, 0x0A, 0x2A, 0x35, 0x18, 0x0B, 0x32, 0x24, 0x55, 0x10, 0x23,
	0x23, 0x3A, 0x28, 0x58, 0x14, 0x20, 0x25, 0x36, 0x07, 0x24, 0x5A, 0x30,
	0x29, 0x2F, 0x0A, 0x59, 0x73, 0x23, 0x36, 0x1C, 0x2C, 0x36, 0x5B, 0x17,
	0x45, 0x0C, 0x7A, 0x3A, 0x16, 0x0F, 0x0E, 0x18, 0x25, 0x55, 0x5E, 0x2D,
	0x2A, 0x55, 0x2B, 0x22, 0x33, 0x17, 0x0A, 0x09, 0x22, 0x0A, 0x30, 0x24,
	0x57, 0x58, 0x5D, 0x69, 0x18, 0x19, 0x1C, 0x44, 0x25, 0x2B, 0x3B, 0x0B,
	0x12, 0x33, 0x2B, 0x14, 0x16, 0x1F, 0x69, 0x3A, 0x08, 0x1B, 0x5E, 0x1A,
	0x19, 0x4E, 0x5A, 0x0D, 0x7B, 0x18, 0x55, 0x2A, 0x22, 0x05, 0x1E, 0x0D,
	0x0B, 0x13, 0x37, 0x09, 0x2B, 0x26, 0x38, 0x13, 0x25, 0x09, 0x37, 0x3E,
	0x3B, 0x58, 0x2A, 0x2D, 0x1A, 0x08, 0x3D, 0x37, 0x3B, 0x39, 0x03, 0x0E,
	0x17, 0x3B, 0x03, 0x20, 0x3B, 0x3B, 0x1E, 0x5A, 0x23, 0x39, 0x15, 0x3C,
	0x12, 0x25, 0x1D, 0x2D, 0x07, 0x29, 0x1A, 0x0E, 0x17, 0x36, 0x31, 0x10,
	0x1F, 0x39, 0x1D, 0x3D, 0x05, 0x15, 0x20, 0x1F, 0x32, 0x37, 0x55, 0x04,
	0x59, 0x2D, 0x70, 0x14, 0x38, 0x56, 0x0D, 0x27, 0x2A, 0x39, 0x18, 0x33,
	0x75, 0x5C, 0x16, 0x5C, 0x1E, 0x3B, 0x3E, 0x2D, 0x39, 0x0E, 0x6D, 0x1A,
	0x17, 0x0A, 0x44, 0x71, 0x47, 0x4E, 0x41, 0x0D, 0x38, 0x47, 0x0B, 0x19,
	0x05, 0x06, 0x1B, 0x54, 0x23, 0x58, 0x12, 0x01, 0x35, 0x23, 0x00, 0x29,
	0x01, 0x51, 0x17, 0x08, 0x34, 0x16, 0x18, 0x0A, 0x3B, 0x01, 0x55, 0x2F,
	0x0A, 0x21, 0x03, 0x07, 0x03, 0x2C, 0x40, 0x27, 0x28, 0x58, 0x02, 0x5B,
	0x69, 0x22, 0x06, 0x21, 0x18, 0x1A, 0x3B, 0x52, 0x27, 0x2E, 0x27, 0x1C,
	0x2E, 0x59, 0x2D, 0x38, 0x01, 0x04, 0x0C, 0x3F, 0x04, 0x04, 0x4A, 0x41,
	0x3C, 0x0B, 0x59, 0x19, 0x5F, 0x2C, 0x71, 0x00, 0x53, 0x3A, 0x1E, 0x1A,
	0x27, 0x31, 0x16, 0x11, 0x7A, 0x1D, 0x10, 0x26, 0x3C, 0x71, 0x36, 0x36,
	0x2A, 0x07, 0x13, 0x43, 0x2C, 0x5D, 0x02, 0x27, 0x47, 0x25, 0x20, 0x13,
	0x6D, 0x22, 0x51, 0x02, 0x38, 0x72, 0x21, 0x0B, 0x0F, 0x3D, 0x2B, 0x43,
	0x06, 0x5B, 0x23, 0x17, 0x5A, 0x2F, 0x1A, 0x0F, 0x2B, 0x0D, 0x58, 0x2A,
	0x1B, 0x34, 0x26, 0x25, 0x29, 0x03, 0x32, 0x36, 0x53, 0x59, 0x52, 0x38,
	0x01, 0x0B, 0x2A, 0x0C, 0x3B, 0x04, 0x33, 0x07, 0x0E, 0x05, 0x2E, 0x19,
	0x1A, 0x11, 0x14, 0x55, 0x26, 0x5C, 0x5C, 0x34, 0x5C, 0x02, 0x26, 0x5C,
	0x25, 0x0F, 0x31, 0x5E, 0x2D, 0x76, 0x38, 0x04, 0x58, 0x40, 0x27, 0x24,
	0x50, 0x5E, 0x3A, 0x29, 0x5E, 0x19, 0x56, 0x0F, 0x75, 0x3B, 0x4E, 0x09,
	0x24, 0x31, 0x15, 0x23, 0x2D, 0x27, 0x08, 0x26, 0x02, 0x22, 0x13, 0x1B,
	0x1E, 0x31, 0x38, 0x11, 0x70, 0x22, 0x2A, 0x39, 0x1C, 0x36, 0x5B, 0x1B,
	0x16, 0x03, 0x0B, 0x1E, 0x0F, 0x0A, 0x1C, 0x7A, 0x26, 0x50, 0x56, 0x5C,
	0x72, 0x0D, 0x31, 0x16, 0x23, 0x76, 0x54, 0x2A, 0x26, 0x05, 0x3B, 0x55,
	0x30, 0x56, 0x3F, 0x04, 0x47, 0x2B, 0x58, 0x08, 0x27, 0x5A, 0x1B, 0x26,
	0x05, 0x70, 0x0F, 0x53, 0x38, 0x5B, 0x77, 0x27, 0x56, 0x39, 0x5E, 0x06,
	0x55, 0x2F, 0x16, 0x01, 0x70, 0x01, 0x31, 0x5D, 0x08, 0x12, 0x5E, 0x53,
	0x2C, 0x12, 0x33, 0x1F, 0x23, 0x5B, 0x40, 0x21, 0x22, 0x0E, 0x19, 0x22,
	0x15, 0x1E, 0x14, 0x07, 0x58, 0x33, 0x2D, 0x0C, 0x19, 0x31, 0x34, 0x0A,
	0x0C, 0x26, 0x11, 0x3B, 0x43, 0x2D, 0x26, 0x03, 0x0F, 0x01, 0x26, 0x5E,
	0x0F, 0x33, 0x20, 0x31, 0x5D, 0x38, 0x06, 0x06, 0x0A, 0x18, 0x00, 0x05,
	0x19, 0x54, 0x41, 0x52, 0x31, 0x20, 0x24, 0x05, 0x27, 0x28, 0x0F, 0x12,
	0x1B, 0x23, 0x23, 0x18, 0x0D, 0x0D, 0x06, 0x11, 0x39, 0x33, 0x08, 0x3C,
	0x77, 0x25, 0x4E, 0x0B, 0x06, 0x17, 0x1E, 0x55, 0x36, 0x39, 0x24, 0x21,
	0x2E, 0x03, 0x0D, 0x26, 0x0B, 0x09, 0x1C, 0x0C, 0x07, 0x15, 0x2A, 0x5A,
	0x3D, 0x1A, 0x2F, 0x32, 0x23, 0x21, 0x2A, 0x54, 0x4E, 0x09, 0x1F, 0x77,
	0x58, 0x55, 0x5C, 0x31, 0x7A, 0x5F, 0x10, 0x26, 0x25, 0x72, 0x55, 0x58,
	0x39, 0x03, 0x0E, 0x2F, 0x58, 0x00, 0x44, 0x37, 0x1C, 0x2E, 0x0F, 0x00,
	0x04, 0x07, 0x51, 0x1F, 0x58, 0x73, 0x55, 0x12, 0x37, 0x39, 0x32, 0x3C,
	0x36, 0x26, 0x5A, 0x76, 0x34, 0x29, 0x2F, 0x04, 0x17, 0x43, 0x05, 0x3D,
	0x3E, 0x15, 0x2E, 0x00, 0x5E, 0x5A, 0x26, 0x5F, 0x32, 0x01, 0x06, 0x30,
	0x2F, 0x50, 0x56, 0x44, 0x34, 0x18, 0x00, 0x1B, 0x11, 0x27, 0x2A, 0x53,
	0x3F, 0x44, 0x74, 0x39, 0x05, 0x24, 0x1B, 0x37, 0x3D, 0x06, 0x3F, 0x03,
	0x70, 0x59, 0x36, 0x14, 0x58, 0x29, 0x19, 0x26, 0x34, 0x0C, 0x11, 0x1F,
	0x2E, 0x3A, 0x3C, 0x37, 0x36, 0x22, 0x2F, 0x39, 0x29, 0x43, 0x50, 0x34,
	0x52, 0x76, 0x22, 0x58, 0x18, 0x32, 0x34, 0x02, 0x59, 0x17, 0x5D, 0x0F,
	0x3B, 0x05, 0x02, 0x44, 0x05, 0x55, 0x26, 0x04, 0x08, 0x31, 0x38, 0x33,
	0x1F, 0x11, 0x72, 0x02, 0x29, 0x3C, 0x19, 0x34, 0x0F, 0x05, 0x41, 0x1E,
	0x76, 0x3B, 0x02, 0x04, 0x22, 0x37, 0x2E, 0x54, 0x5D, 0x12, 0x77, 0x00,
	0x30, 0x3B, 0x3D, 0x20, 0x3A, 0x55, 0x36, 0x0E, 0x71, 0x2F, 0x51, 0x0F,
	0x2D, 0x29, 0x36, 0x24, 0x28, 0x06, 0x38, 0x5C, 0x31, 0x00, 0x38, 0x34,
	0x1B, 0x03, 0x5F, 0x5D, 0x23, 0x15, 0x59, 0x39, 0x31, 0x16, 0x36, 0x00,
	0x3C, 0x12, 0x38, 0x3E, 0x2E, 0x1C, 0x1E, 0x37, 0x1E, 0x4E, 0x58, 0x27,
	0x7B, 0x35, 0x4A, 0x08, 0x23, 0x28, 0x1D, 0x09, 0x23, 0x5B, 0x0D, 0x34,
	0x2E, 0x26, 0x02, 0x01, 0x06, 0x29, 0x04, 0x0F, 0x0D, 0x47, 0x29, 0x1F,
	0x28, 0x2D, 0x19, 0x09, 0x01, 0x5D, 0x1B, 0x3C, 0x22, 0x3D, 0x38, 0x29,
	0x03, 0x57, 0x04, 0x02, 0x77, 0x20, 0x06, 0x2A, 0x26, 0x71, 0x39, 0x52,
	0x36, 0x27, 0x2A, 0x3E, 0x36, 0x39, 0x53, 0x04, 0x07, 0x36, 0x2C, 0x5C,
	0x1B, 0x26, 0x11, 0x0F, 0x52, 0x36, 0x39, 0x14, 0x56, 0x3A, 0x04, 0x1D,
	0x34, 0x59, 0x09, 0x77, 0x1D, 0x23, 0x3E, 0x3E, 0x30, 0x06, 0x02, 0x0C,
	0x5A, 0x01, 0x19, 0x22, 0x1A, 0x3B, 0x18, 0x24, 0x35, 0x1C, 0x38, 0x69,
	0x1A, 0x59, 0x07, 0x27, 0x05, 0x26, 0x4E, 0x19, 0x12, 0x2E, 0x3F, 0x1B,
	0x3E, 0x20, 0x20, 0x34, 0x57, 0x16, 0x58, 0x77, 0x06, 0x0F, 0x45, 0x5E,
	0x0E, 0x05, 0x23, 0x39, 0x1E, 0x16, 0x5E, 0x56, 0x1F, 0x58, 0x1A, 0x01,
	0x53, 0x16, 0x20, 0x20, 0x47, 0x2B, 0x17, 0x21, 0x23, 0x1F, 0x24, 0x41,
	0x02, 0x03, 0x20, 0x15, 0x2D, 0x52, 0x0F, 0x3C, 0x0E, 0x16, 0x09, 0x28,
	0x3E, 0x13, 0x01, 0x26, 0x34, 0x47, 0x25, 0x5C, 0x1F, 0x25, 0x08, 0x09,
	0x0B, 0x26, 0x30, 0x5B, 0x58, 0x37, 0x0D, 0x31, 0x5D, 0x32, 0x1D, 0x3C,
	0x2E, 0x5C, 0x37, 0x23, 0x26, 0x2B, 0x5A, 0x3B, 0x3F, 0x3F, 0x16, 0x54,
	0x04, 0x45, 0x2D, 0x74, 0x04, 0x1B, 0x1B, 0x29, 0x17, 0x1B, 0x4A, 0x01,
	0x1B, 0x13, 0x58, 0x18, 0x58, 0x0D, 0x69, 0x2B, 0x32, 0x29, 0x5D, 0x21,
	0x43, 0x03, 0x14, 0x3E, 0x71, 0x5E, 0x0B, 0x45, 0x5E, 0x69, 0x05, 0x2B,
	0x0C, 0x01, 0x0D, 0x16, 0x29, 0x2F, 0x06, 0x24, 0x59, 0x0F, 0x02, 0x1F,
	0x1A, 0x05, 0x4A, 0x59, 0x52, 0x05, 0x5F, 0x56, 0x0C, 0x00, 0x34, 0x06,
	0x15, 0x45, 0x2E, 0x16, 0x05, 0x34, 0x39, 0x1F, 0x08, 0x1B, 0x50, 0x5B,
	0x04, 0x23, 0x02, 0x56, 0x0C, 0x0D, 0x15, 0x0B, 0x18, 0x07, 0x1E, 0x34,
	0x5D, 0x0B, 0x56, 0x00, 0x09, 0x04, 0x10, 0x57, 0x01, 0x71, 0x18, 0x52,
	0x41, 0x5F, 0x69, 0x55, 0x23, 0x39, 0x5F, 0x24, 0x24, 0x0C, 0x58, 0x5A,
	0x77, 0x04, 0x2C, 0x22, 0x40, 0x2F, 0x43, 0x2A, 0x59, 0x19, 0x06, 0x5C,
	0x59, 0x0C, 0x19, 0x27, 0x2A, 0x1B, 0x34, 0x23, 0x71, 0x02, 0x2C, 0x0D,
	0x38, 0x27, 0x14, 0x56, 0x0B, 0x5D, 0x36, 0x05, 0x56, 0x5C, 0x2D, 0x38,
	0x29, 0x59, 0x1A, 0x01, 0x04, 0x39, 0x55, 0x5D, 0x3B, 0x09, 0x54, 0x35,
	0x5A, 0x39, 0x04, 0x38, 0x50, 0x56, 0x58, 0x20, 0x5F, 0x07, 0x2C, 0x18,
	0x76, 0x5D, 0x29, 0x3A, 0x3D, 0x33, 0x5B, 0x33, 0x0C, 0x3E, 0x31, 0x07,
	0x53, 0x16, 0x0A, 0x0A, 0x06, 0x53, 0x16, 0x58, 0x6D, 0x0F, 0x22, 0x2F,
	0x21, 0x23, 0x00, 0x57, 0x1B, 0x32, 0x0A, 0x1C, 0x09, 0x20, 0x0A, 0x37,
	0x04, 0x02, 0x03, 0x06, 0x75, 0x5E, 0x05, 0x5F, 0x11, 0x00, 0x0B, 0x4E,
	0x5F, 0x0A, 0x01, 0x20, 0x04, 0x3C, 0x05, 0x2A, 0x5E, 0x32, 0x2D, 0x5C,
	0x26, 0x35, 0x02, 0x1B, 0x33, 0x14, 0x5F, 0x00, 0x5C, 0x06, 0x7B, 0x0A,
	0x24, 0x57, 0x3B, 0x13, 0x02, 0x20, 0x06, 0x19, 0x29, 0x1C, 0x02, 0x56,
	0x38, 0x30, 0x22, 0x39, 0x14, 0x1E, 0x1B, 0x0A, 0x13, 0x36, 0x3B, 0x71,
	0x20, 0x23, 0x1E, 0x2E, 0x30, 0x2B, 0x14, 0x1E, 0x0F, 0x20, 0x16, 0x4E,
	0x5B, 0x3B, 0x75, 0x3F, 0x18, 0x2C, 0x5D, 0x70, 0x23, 0x16, 0x0B, 0x5C,
	0x0A, 0x05, 0x3B, 0x21, 0x2C, 0x33, 0x43, 0x4A, 0x08, 0x1D, 0x1A, 0x3F,
	0x35, 0x1E, 0x52, 0x34, 0x28, 0x4E, 0x0D, 0x22, 0x75, 0x43, 0x0C, 0x37,
	0x2E, 0x34, 0x1F, 0x08, 0x57, 0x2E, 0x21, 0x26, 0x4E, 0x2C, 0x5C, 0x71,
	0x5F, 0x02, 0x5F, 0x09, 0x18, 0x55, 0x39, 0x23, 0x25, 0x08, 0x1C, 0x55,
	0x45, 0x09, 0x0E, 0x5F, 0x0A, 0x1A, 0x32, 0x06, 0x3A, 0x52, 0x3C, 0x5F,
	0x23, 0x02, 0x39, 0x28, 0x44, 0x36, 0x5B, 0x18, 0x36, 0x3E, 0x10, 0x25,
	0x11, 0x56, 0x5A, 0x71, 0x20, 0x06, 0x57, 0x33, 0x04, 0x54, 0x52, 0x21,
	0x24, 0x34, 0x20, 0x35, 0x34, 0x05, 0x17, 0x28, 0x0E, 0x01, 0x01, 0x29,
	0x20, 0x3B, 0x1E, 0x59, 0x7B, 0x0F, 0x08, 0x26, 0x2F, 0x76, 0x5D, 0x52,
	0x04, 0x26, 0x29, 0x5A, 0x51, 0x5A, 0x08, 0x0B, 0x03, 0x30, 0x1E, 0x27,
	0x1A, 0x54, 0x51, 0x0D, 0x1F, 0x37, 0x3A, 0x05, 0x56, 0x44, 0x38, 0x0E,
	0x0B, 0x0A, 0x5A, 0x09, 0x05, 0x20, 0x34, 0x00, 0x1B, 0x1A, 0x0F, 0x59,
	0x3B, 0x2B, 0x0F, 0x13, 0x0A, 0x5E, 0x35, 0x43, 0x4A, 0x07, 0x12, 0x35,
	0x1E, 0x35, 0x58, 0x13, 0x3B, 0x2B, 0x50, 0x56, 0x32, 0x06, 0x1E, 0x4E,
	0x06, 0x58, 0x1A, 0x54, 0x51, 0x34, 0x58, 0x77, 0x27, 0x1B, 0x0C, 0x58,
	0x08, 0x00, 0x18, 0x23, 0x3C, 0x77, 0x1A, 0x0F, 0x59, 0x24, 0x2C, 0x47,
	0x18, 0x0F, 0x3D, 0x0E, 0x0B, 0x0C, 0x2F, 0x1A, 0x0E, 0x59, 0x4E, 0x3F,
	0x06, 0x2A, 0x0E, 0x36, 0x56, 0x25, 0x32, 0x0F, 0x18, 0x56, 0x33, 0x0A,
	0x3B, 0x13, 0x00, 0x3C, 0x06, 0x5B, 0x4A, 0x01, 0x38, 0x27, 0x06, 0x38,
	0x1C, 0x3D, 0x31, 0x07, 0x57, 0x28, 0x1A, 0x77, 0x0A, 0x50, 0x08, 0x38,
	0x37, 0x0F, 0x15, 0x24, 0x13, 0x71, 0x5E, 0x2B, 0x5E, 0x53, 0x75, 0x04,
	0x4A, 0x5F, 0x1D, 0x71, 0x3F, 0x0A, 0x1E, 0x5C, 0x21, 0x02, 0x32, 0x07,
	0x58, 0x30, 0x2B, 0x14, 0x3D, 0x5F, 0x28, 0x3F, 0x22, 0x34, 0x08, 0x6D,
	0x04, 0x33, 0x39, 0x3B, 0x24, 0x43, 0x33, 0x58, 0x12, 0x13, 0x34, 0x2F,
	0x2F, 0x0A, 0x31, 0x26, 0x0E, 0x1A, 0x21, 0x01, 0x0E, 0x4E, 0x18, 0x11,
	0x2A, 0x0E, 0x27, 0x3C, 0x1F, 0x2A, 0x23, 0x2E, 0x45, 0x3C, 0x75, 0x3E,
	0x05, 0x17, 0x24, 0x11, 0x5B, 0x2C, 0x59, 0x0E, 0x28, 0x15, 0x4E, 0x0A,
	0x40, 0x75, 0x02, 0x2D, 0x0F, 0x1E, 0x24, 0x47, 0x34, 0x0C, 0x25, 0x2C,
	0x29, 0x58, 0x5B, 0x0D, 0x3B, 0x3A, 0x15, 0x04, 0x40, 0x16, 0x0E, 0x25,
	0x24, 0x0C, 0x1A, 0x5A, 0x03, 0x18, 0x5C, 0x21, 0x47, 0x32, 0x21, 0x03,
	0x26, 0x5F, 0x2F, 0x41, 0x1E, 0x7B, 0x58, 0x58, 0x03, 0x1D, 0x29, 0x5D,
	0x31, 0x28, 0x0D, 0x12, 0x1F, 0x31, 0x56, 0x5F, 0x18, 0x15, 0x28, 0x01,
	0x21, 0x01, 0x5F, 0x0B, 0x3F, 0x08, 0x01, 0x55, 0x17, 0x41, 0x1B, 0x74,
	0x2B, 0x0B, 0x38, 0x5F, 0x23, 0x16, 0x57, 0x34, 0x02, 0x0A, 0x00, 0x18,
	0x5B, 0x1D, 0x3A, 0x2D, 0x12, 0x41, 0x5D, 0x27, 0x2B, 0x4A, 0x0D, 0x5A,
	0x34, 0x20, 0x11, 0x06, 0x53, 0x06, 0x3C, 0x08, 0x38, 0x1E, 0x6D, 0x55,
	0x56, 0x1A, 0x0F, 0x38, 0x47, 0x54, 0x17, 0x5B, 0x0A, 0x0E, 0x52, 0x45,
	0x3E, 0x17, 0x2F, 0x13, 0x04, 0x00, 0x10, 0x03, 0x4E, 0x1D, 0x32, 0x05,
	0x55, 0x03, 0x41, 0x32, 0x28, 0x08, 0x54, 0x5F, 0x08, 0x72, 0x2B, 0x34,
	0x5C, 0x0D, 0x0F, 0x14, 0x19, 0x2A, 0x24, 0x06, 0x3B, 0x16, 0x18, 0x05,
	0x24, 0x08, 0x13, 0x0A, 0x1D, 0x05, 0x5F, 0x25, 0x00, 0x11, 0x34, 0x0E,
	0x31, 0x1C, 0x1B, 0x0C, 0x1A, 0x25, 0x5D, 0x0E, 0x28, 0x06, 0x05, 0x19,
	0x13, 0x0C, 0x14, 0x2F, 0x36, 0x31, 0x08, 0x5B, 0x2F, 0x06, 0x03, 0x27,
	0x5E, 0x3B, 0x5B, 0x22, 0x0A, 0x08, 0x0C, 0x1E, 0x18, 0x0C, 0x21, 0x50,
	0x5B, 0x5E, 0x23, 0x38, 0x07, 0x27, 0x22, 0x15, 0x20, 0x0F, 0x09, 0x40,
	0x2E, 0x26, 0x09, 0x58, 0x58, 0x23, 0x5F, 0x4A, 0x19, 0x39, 0x38, 0x18,
	0x2F, 0x05, 0x3D, 0x0C, 0x3A, 0x4E, 0x58, 0x52, 0x30, 0x47, 0x20, 0x07,
	0x5F, 0x1A, 0x0B, 0x59, 0x56, 0x3D, 0x2C, 0x3B, 0x27, 0x5D, 0x2D, 0x07,
	0x39, 0x04, 0x38, 0x03, 0x3A, 0x15, 0x14, 0x3E, 0x3C, 0x3A, 0x21, 0x35,
	0x1B, 0x58, 0x30, 0x29, 0x0C, 0x39, 0x38, 0x0C, 0x09, 0x39, 0x05, 0x13,
	0x23, 0x0E, 0x15, 0x58, 0x1D, 0x14, 0x35, 0x11, 0x3C, 0x2D, 0x3B, 0x1A,
	0x32, 0x5C, 0x26, 0x05, 0x04, 0x13, 0x0A, 0x18, 0x32, 0x47, 0x2F, 0x04,
	0x5F, 0x14, 0x5E, 0x53, 0x57, 0x01, 0x2B, 0x3E, 0x29, 0x08, 0x01, 0x03,
	0x35, 0x31, 0x2B, 0x53, 0x1B, 0x3A, 0x4A, 0x20, 0x0C, 0x07, 0x16, 0x13,
	0x0F, 0x25, 0x72, 0x3B, 0x23, 0x29, 0x44, 0x04, 0x1E, 0x30, 0x1B, 0x1E,
	0x0B, 0x14, 0x58, 0x36, 0x0E, 0x34, 0x3C, 0x0C, 0x0C, 0x05, 0x27, 0x09,
	0x28, 0x3D, 0x32, 0x09, 0x09, 0x50, 0x5D, 0x59, 0x01, 0x3A, 0x54, 0x1D,
	0x44, 0x33, 0x26, 0x31, 0x19, 0x05, 0x06, 0x14, 0x59, 0x0A, 0x0D, 0x75,
	0x05, 0x25, 0x3B, 0x1D, 0x08, 0x15, 0x38, 0x0C, 0x27, 0x69, 0x43, 0x0A,
	0x5A, 0x2F, 0x13, 0x5E, 0x57, 0x36, 0x09, 0x38, 0x54, 0x2C, 0x0F, 0x2E,
	0x21, 0x22, 0x20, 0x04, 0x05, 0x35, 0x04, 0x15, 0x0A, 0x52, 0x21, 0x43,
	0x0D, 0x00, 0x1E, 0x0A, 0x3C, 0x56, 0x2F, 0x0E, 0x13, 0x28, 0x1B, 0x5C,
	0x26, 0x0D, 0x18, 0x39, 0x08, 0x23, 0x0E, 0x23, 0x14, 0x3B, 0x0E, 0x16,
	0x01, 0x57, 0x16, 0x1D, 0x0F, 0x3B, 0x16, 0x22, 0x32, 0x1A, 0x38, 0x18,
	0x5D, 0x38, 0x26, 0x43, 0x51, 0x0C, 0x0E, 0x75, 0x43, 0x20, 0x57, 0x59,
	0x73, 0x1F, 0x38, 0x00, 0x2F, 0x1B, 0x00, 0x2D, 0x5D, 0x11, 0x31, 0x58,
	0x59, 0x04, 0x21, 0x71, 0x01, 0x4A, 0x5B, 0x52, 0x70, 0x43, 0x39, 0x04,
	0x07, 0x27, 0x54, 0x09, 0x3C, 0x20, 0x7B, 0x3E, 0x31, 0x14, 0x1C, 0x27,
	0x04, 0x19, 0x3C, 0x2D, 0x30, 0x5A, 0x17, 0x3B, 0x0E, 0x10, 0x43, 0x30,
	0x18, 0x32, 0x25, 0x25, 0x50, 0x29, 0x44, 0x18, 0x5F, 0x08, 0x07, 0x01,
	0x23, 0x23, 0x4E, 0x09, 0x12, 0x77, 0x35, 0x56, 0x2C, 0x33, 0x07, 0x5A,
	0x19, 0x20, 0x5A, 0x38, 0x28, 0x1B, 0x20, 0x28, 0x74, 0x16, 0x05, 0x0D,
	0x19, 0x38, 0x2A, 0x2F, 0x56, 0x1E, 0x28, 0x47, 0x35, 0x5D, 0x40, 0x2B,
	0x5F, 0x19, 0x45, 0x39, 0x04, 0x59, 0x57, 0x29, 0x52, 0x1B, 0x5F, 0x30,
	0x5C, 0x1E, 0x00, 0x1A, 0x05, 0x1F, 0x1F, 0x2C, 0x24, 0x17, 0x28, 0x21,
	0x70, 0x23, 0x19, 0x3F, 0x53, 0x04, 0x2D, 0x0F, 0x3C, 0x44, 0x05, 0x20,
	0x12, 0x16, 0x0E, 0x24, 0x18, 0x0D, 0x2B, 0x01, 0x12, 0x05, 0x00, 0x5E,
	0x12, 0x2C, 0x0B, 0x51, 0x3C, 0x59, 0x12, 0x05, 0x17, 0x1D, 0x0D, 0x17,
	0x00, 0x20, 0x0D, 0x0F, 0x12, 0x2D, 0x0A, 0x26, 0x52, 0x74, 0x38, 0x06,
	0x21, 0x5B, 0x76, 0x47, 0x0D, 0x07, 0x44, 0x34, 0x38, 0x0F, 0x09, 0x40,
	0x21, 0x3C, 0x30, 0x56, 0x0C, 0x25, 0x16, 0x33, 0x22, 0x2C, 0x28, 0x05,
	0x07, 0x39, 0x58, 0x06, 0x2B, 0x15, 0x3E, 0x53, 0x25, 0x0B, 0x4E, 0x20,
	0x1D, 0x3A, 0x2A, 0x0B, 0x0D, 0x59, 0x0D, 0x5D, 0x2B, 0x2B, 0x06, 0x12,
	0x5A, 0x4E, 0x3B, 0x5D, 0x26, 0x55, 0x33, 0x1F, 0x5A, 0x69, 0x16, 0x14,
	0x16, 0x3B, 0x09, 0x08, 0x0E, 0x5D, 0x38, 0x2F, 0x43, 0x33, 0x05, 0x52,
	0x23, 0x54, 0x0F, 0x06, 0x11, 0x77, 0x1F, 0x32, 0x3E, 0x00, 0x76, 0x06,
	0x05, 0x25, 0x12, 0x23, 0x5D, 0x51, 0x1A, 0x1F, 0x37, 0x5F, 0x12, 0x1C,
	0x5E, 0x20, 0x06, 0x0B, 0x1A, 0x07, 0x37, 0x02, 0x32, 0x05, 0x20, 0x28,
	0x05, 0x52, 0x5D, 0x28, 0x25, 0x54, 0x4A, 0x5B, 0x1D, 0x23, 0x3C, 0x2F,
	0x22, 0x5E, 0x38, 0x5C, 0x2F, 0x0B, 0x1F, 0x0F, 0x09, 0x23, 0x41, 0x1F,
	0x21, 0x3B, 0x22, 0x09, 0x5B, 0x77, 0x0F, 0x29, 0x36, 0x5E, 0x76, 0x09,
	0x56, 0x0C, 0x2D, 0x29, 0x16, 0x39, 0x07, 0x02, 0x11, 0x08, 0x00, 0x34,
	0x1F, 0x09, 0x2A, 0x29, 0x06, 0x02, 0x71, 0x0E, 0x4A, 0x3D, 0x2A, 0x30,
	0x07, 0x2C, 0x1F, 0x52, 0x16, 0x59, 0x35, 0x01, 0x5C, 0x36, 0x0A, 0x34,
	0x29, 0x09, 0x2F, 0x3B, 0x18, 0x1C, 0x33, 0x16, 0x21, 0x19, 0x1E, 0x58,
	0x35, 0x59, 0x3B, 0x37, 0x2E, 0x30, 0x04, 0x19, 0x1D, 0x07, 0x74, 0x43,
	0x04, 0x39, 0x1B, 0x18, 0x34, 0x38, 0x3E, 0x06, 0x30, 0x1C, 0x06, 0x14,
	0x05, 0x0A, 0x2E, 0x07, 0x5E, 0x33, 0x38, 0x08, 0x53, 0x0A, 0x0E, 0x75,
	0x3C, 0x02, 0x20, 0x5A, 0x14, 0x06, 0x11, 0x3E, 0x0F, 0x20, 0x1C, 0x2A,
	0x2A, 0x21, 0x2D, 0x58, 0x4A, 0x58, 0x39, 0x18, 0x59, 0x15, 0x17, 0x1B,
	0x13, 0x14, 0x4A, 0x1B, 0x3D, 0x25, 0x1F, 0x4E, 0x5C, 0x22, 0x1B, 0x58,
	0x3B, 0x24, 0x05, 0x18, 0x58, 0x4A, 0x00, 0x2D, 0x76, 0x0E, 0x38, 0x20,
	0x22, 0x31, 0x54, 0x04, 0x1A, 0x1F, 0x76, 0x15, 0x09, 0x23, 0x02, 0x2D,
	0x0E, 0x29, 0x2D, 0x06, 0x7B, 0x36, 0x30, 0x03, 0x11, 0x29, 0x5E, 0x02,
	0x5D, 0x2F, 0x7A, 0x5A, 0x0C, 0x1E, 0x5B, 0x2A, 0x0A, 0x23, 0x1B, 0x0F,
	0x10, 0x19, 0x24, 0x08, 0x0C, 0x25, 0x58, 0x3B, 0x3B, 0x2D, 0x0D, 0x47,
	0x29, 0x22, 0x01, 0x0B, 0x25, 0x57, 0x59, 0x58, 0x13, 0x43, 0x14, 0x08,
	0x1D, 0x76, 0x5F, 0x3B, 0x0B, 0x06, 0x05, 0x54, 0x58, 0x0D, 0x5D, 0x71,
	0x5E, 0x0E, 0x00, 0x2E, 0x69, 0x38, 0x32, 0x36, 0x5A, 0x76, 0x54, 0x10,
	0x57, 0x5D, 0x35, 0x58, 0x15, 0x07, 0x1A, 0x38, 0x3D, 0x2E, 0x24, 0x44,
	0x29, 0x28, 0x0B, 0x01, 0x0D, 0x27, 0x14, 0x25, 0x3A, 0x1A, 0x0C, 0x18,
	0x55, 0x1B, 0x52, 0x0A, 0x05, 0x09, 0x25, 0x24, 0x05, 0x28, 0x30, 0x02,
	0x1F, 0x34, 0x3D, 0x3B, 0x59, 0x1F, 0x00, 0x1C, 0x32, 0x0F, 0x1E, 0x6D,
	0x55, 0x16, 0x17, 0x5C, 0x10, 0x23, 0x57, 0x37, 0x2E, 0x72, 0x01, 0x38,
	0x38, 0x38, 0x76, 0x35, 0x57, 0x14, 0x09, 0x69, 0x47, 0x02, 0x1A, 0x05,
	0x2E, 0x5A, 0x05, 0x3F, 0x40, 0x16, 0x18, 0x53, 0x2B, 0x2A, 0x71, 0x02,
	0x4E, 0x0D, 0x11, 0x10, 0x3C, 0x08, 0x41, 0x26, 0x07, 0x2E, 0x56, 0x1E,
	0x0D, 0x01, 0x2D, 0x4A, 0x5D, 0x31, 0x2A, 0x35, 0x2F, 0x25, 0x27, 0x2C,
	0x47, 0x57, 0x02, 0x23, 0x01, 0x03, 0x2C, 0x08, 0x31, 0x3A, 0x5B, 0x00,
	0x5B, 0x28, 0x33, 0x25, 0x28, 0x23, 0x09, 0x70, 0x02, 0x07, 0x00, 0x2C,
	0x7B, 0x00, 0x2F, 0x19, 0x44, 0x0C, 0x5E, 0x54, 0x29, 0x38, 0x70, 0x28,
	0x38, 0x5A, 0x1E, 0x08, 0x02, 0x20, 0x3B, 0x27, 0x35, 0x59, 0x15, 0x08,
	0x05, 0x77, 0x23, 0x58, 0x08, 0x1F, 0x13, 0x0D, 0x55, 0x0B, 0x32, 0x24,
	0x09, 0x12, 0x3D, 0x3C, 0x0A, 0x5E, 0x31, 0x39, 0x58, 0x38, 0x47, 0x52,
	0x01, 0x53, 0x0E, 0x07, 0x54, 0x06, 0x12, 0x30, 0x15, 0x23, 0x5A, 0x28,
	0x0B, 0x1A, 0x13, 0x26, 0x5C, 0x24, 0x25, 0x23, 0x29, 0x04, 0x7B, 0x21,
	0x33, 0x2C, 0x0F, 0x71, 0x5E, 0x29, 0x56, 0x20, 0x15, 0x29, 0x37, 0x56,
	0x44, 0x38, 0x2B, 0x50, 0x5A, 0x2E, 0x36, 0x21, 0x35, 0x1B, 0x19, 0x37,
	0x2F, 0x3B, 0x1A, 0x09, 0x75, 0x05, 0x56, 0x3C, 0x22, 0x12, 0x0E, 0x59,
	0x3D, 0x24, 0x2C, 0x55, 0x04, 0x0F, 0x3F, 0x17, 0x5B, 0x57, 0x05, 0x5F,
	0x75, 0x55, 0x26, 0x3A, 0x44, 0x28, 0x5B, 0x24, 0x5A, 0x23, 0x72, 0x02,
	0x37, 0x04, 0x18, 0x37, 0x5A, 0x39, 0x5E, 0x19, 0x26, 0x1F, 0x18, 0x05,
	0x1A, 0x0C, 0x0E, 0x32, 0x3C, 0x3A, 0x11, 0x5D, 0x07, 0x0B, 0x05, 0x10,
	0x2A, 0x02, 0x3C, 0x09, 0x2C, 0x3B, 0x37, 0x2C, 0x5C, 0x6D, 0x0A, 0x2C,
	0x03, 0x5F, 0x11, 0x25, 0x30, 0x59, 0x2D, 0x6D, 0x36, 0x2E, 0x05, 0x0E,
	0x70, 0x24, 0x25, 0x58, 0x01, 0x77, 0x34, 0x53, 0x3D, 0x33, 0x37, 0x27,
	0x39, 0x27, 0x01, 0x71, 0x5F, 0x19, 0x45, 0x2D, 0x38, 0x55, 0x09, 0x05,
	0x24, 0x28, 0x0E, 0x23, 0x18, 0x40, 0x27, 0x0A, 0x06, 0x17, 0x44, 0x2E,
	0x29, 0x26, 0x00, 0x0D, 0x75, 0x5B, 0x1B, 0x01, 0x18, 0x01, 0x14, 0x57,
	0x45, 0x09, 0x2B, 0x3B, 0x23, 0x01, 0x07, 0x0A, 0x08, 0x2F, 0x5A, 0x3F,
	0x7A, 0x38, 0x52, 0x39, 0x24, 0x76, 0x14, 0x3B, 0x0B, 0x33, 0x12, 0x3A,
	0x19, 0x18, 0x3A, 0x73, 0x14, 0x23, 0x59, 0x27, 0x0E, 0x02, 0x23, 0x2C,
	0x3D, 0x07, 0x5A, 0x28, 0x57, 0x29, 0x30, 0x1D, 0x2D, 0x17, 0x5B, 0x38,
	0x26, 0x06, 0x0A, 0x27, 0x6D, 0x05, 0x35, 0x29, 0x09, 0x25, 0x1B, 0x59,
	0x23, 0x2F, 0x10, 0x03, 0x51, 0x0F, 0x11, 0x06, 0x04, 0x19, 0x37, 0x08,
	0x2F, 0x23, 0x0B, 0x41, 0x03, 0x0A, 0x04, 0x15, 0x21, 0x5D, 0x10, 0x20,
	0x51, 0x3C, 0x2A, 0x72, 0x58, 0x14, 0x18, 0x1C, 0x18, 0x3D, 0x12, 0x18,
	0x05, 0x0D, 0x5D, 0x20, 0x1C, 0x29, 0x7B, 0x47, 0x4A, 0x03, 0x02, 0x06,
	0x2B, 0x00, 0x38, 0x52, 0x26, 0x1A, 0x39, 0x3C, 0x11, 0x06, 0x5B, 0x0C,
	0x3E, 0x1B, 0x33, 0x25, 0x14, 0x28, 0x19, 0x74, 0x09, 0x04, 0x28, 0x2C,
	0x24, 0x1D, 0x34, 0x38, 0x33, 0x38, 0x18, 0x17, 0x5F, 0x53, 0x15, 0x0E,
	0x19, 0x24, 0x3E, 0x6D, 0x38, 0x03, 0x1F, 0x03, 0x73, 0x2E, 0x03, 0x14,
	0x06, 0x37, 0x14, 0x35, 0x36, 0x44, 0x14, 0x19, 0x37, 0x3A, 0x1D, 0x2B,
	0x55, 0x2B, 0x01, 0x3C, 0x24, 0x1D, 0x34, 0x58, 0x40, 0x14, 0x47, 0x39,
	0x5C, 0x3C, 0x2B, 0x09, 0x56, 0x06, 0x28, 0x1B, 0x3D, 0x03, 0x07, 0x2E,
	0x12, 0x2E, 0x16, 0x09, 0x06, 0x16, 0x5B, 0x1B, 0x07, 0x40, 0x18, 0x02,
	0x29, 0x5B, 0x0F, 0x7B, 0x15, 0x59, 0x56, 0x3F, 0x2A, 0x09, 0x59, 0x5C,
	0x24, 0x0F, 0x0A, 0x15, 0x39, 0x3B, 0x2A, 0x18, 0x50, 0x39, 0x20, 0x20,
	0x14, 0x55, 0x5F, 0x3C, 0x36, 0x15, 0x2D, 0x21, 0x1D, 0x69, 0x59, 0x52,
	0x08, 0x22, 0x3A, 0x00, 0x00, 0x0A, 0x08, 0x18, 0x36, 0x2B, 0x0D, 0x3D,
	0x6D, 0x3B, 0x02, 0x05, 0x2E, 0x26, 0x58, 0x17, 0x20, 0x40, 0x73, 0x19,
	0x18, 0x3D, 0x53, 0x77, 0x5C, 0x02, 0x26, 0x52, 0x74, 0x25, 0x0C, 0x5D,
	0x2C, 0x76, 0x54, 0x32, 0x14, 0x12, 0x7A, 0x2B, 0x39, 0x3A, 0x21, 0x37,
	0x39, 0x05, 0x14, 0x02, 0x77, 0x47, 0x30, 0x57, 0x2A, 0x77, 0x5F, 0x2E,
	0x20, 0x02, 0x12, 0x0D, 0x0F, 0x28, 0x03, 0x77, 0x35, 0x12, 0x26, 0x1A,
	0x12, 0x0B, 0x58, 0x26, 0x19, 0x3A, 0x1F, 0x59, 0x38, 0x22, 0x0D, 0x27,
	0x2B, 0x3A, 0x09, 0x37, 0x54, 0x07, 0x41, 0x40, 0x13, 0x5B, 0x58, 0x17,
	0x59, 0x26, 0x20, 0x54, 0x29, 0x0C, 0x70, 0x23, 0x34, 0x36, 0x1E, 0x08,
	0x3A, 0x4A, 0x45, 0x2F, 0x00, 0x03, 0x10, 0x5E, 0x3B, 0x75, 0x3D, 0x57,
	0x5C, 0x2C, 0x09, 0x2F, 0x52, 0x09, 0x2F, 0x38, 0x3E, 0x12, 0x3D, 0x0C,
	0x36, 0x43, 0x02, 0x58, 0x09, 0x18, 0x43, 0x57, 0x57, 0x05, 0x2F, 0x5A,
	0x54, 0x0B, 0x1A, 0x25, 0x08, 0x51, 0x36, 0x52, 0x01, 0x21, 0x4E, 0x25,
	0x44, 0x36, 0x38, 0x10, 0x28, 0x3B, 0x77, 0x06, 0x30, 0x56, 0x06, 0x0F,
	0x01, 0x28, 0x5F, 0x11, 0x0C, 0x14, 0x29, 0x1A, 0x2C, 0x38, 0x39, 0x50,
	0x0C, 0x40, 0x12, 0x36, 0x38, 0x1E, 0x0A, 0x0D, 0x3E, 0x11, 0x0A, 0x09,
	0x0F, 0x43, 0x55, 0x17, 0x22, 0x0E, 0x35, 0x15, 0x14, 0x05, 0x31, 0x1D,
	0x14, 0x3D, 0x11, 0x37, 0x22, 0x2F, 0x5D, 0x5C, 0x74, 0x22, 0x16, 0x5D,
	0x2E, 0x76, 0x38, 0x24, 0x17, 0x0C, 0x0F, 0x47, 0x27, 0x18, 0x33, 0x7A,
	0x43, 0x19, 0x5A, 0x05, 0x23, 0x08, 0x2A, 0x02, 0x1A, 0x73, 0x5D, 0x02,
	0x27, 0x31, 0x05, 0x0A, 0x27, 0x0B, 0x2A, 0x76, 0x0D, 0x04, 0x0C, 0x59,
	0x71, 0x0B, 0x59, 0x5D, 0x3E, 0x00, 0x22, 0x17, 0x57, 0x1F, 0x13, 0x01,
	0x25, 0x23, 0x1F, 0x77, 0x02, 0x0E, 0x3E, 0x38, 0x0E, 0x3E, 0x56, 0x0B,
	0x33, 0x37, 0x16, 0x19, 0x56, 0x24, 0x08, 0x21, 0x31, 0x58, 0x20, 0x00,
	0x0A, 0x14, 0x24, 0x07, 0x28, 0x5B, 0x2D, 0x07, 0x59, 0x73, 0x0F, 0x2E,
	0x36, 0x2C, 0x32, 0x59, 0x28, 0x00, 0x5B, 0x32, 0x0F, 0x00, 0x1F, 0x3A,
	0x72, 0x2B, 0x0B, 0x18, 0x0F, 0x34, 0x1E, 0x3B, 0x05, 0x32, 0x17, 0x3C,
	0x09, 0x2F, 0x24, 0x73, 0x27, 0x2E, 0x24, 0x05, 0x6D, 0x34, 0x27, 0x26,
	0x1F, 0x7A, 0x58, 0x14, 0x14, 0x33, 0x26, 0x2F, 0x15, 0x16, 0x52, 0x2C,
	0x02, 0x29, 0x2F, 0x05, 0x6D, 0x1C, 0x55, 0x08, 0x58, 0x11, 0x3A, 0x0C,
	0x1B, 0x5D, 0x16, 0x21, 0x10, 0x59, 0x39, 0x10, 0x06, 0x31, 0x26, 0x0E,
	0x1A, 0x2B, 0x2B, 0x2A, 0x52, 0x7B, 0x5E, 0x00, 0x5D, 0x39, 0x77, 0x21,
	0x0C, 0x16, 0x2A, 0x2A, 0x19, 0x05, 0x2B, 0x5A, 0x76, 0x1A, 0x0D, 0x00,
	0x32, 0x30, 0x1E, 0x26, 0x1E, 0x3A, 0x2F, 0x09, 0x23, 0x1B, 0x33, 0x00,
	0x06, 0x0A, 0x0D, 0x38, 0x0E, 0x0E, 0x3B, 0x5D, 0x5C, 0x07, 0x36, 0x51,
	0x56, 0x25, 0x04, 0x59, 0x53, 0x23, 0x03, 0x76, 0x3E, 0x11, 0x18, 0x2F,
	0x28, 0x03, 0x05, 0x0B, 0x19, 0x2C, 0x27, 0x3B, 0x3D, 0x1F, 0x6D, 0x43,
	0x59, 0x39, 0x27, 0x26, 0x3A, 0x37, 0x21, 0x5D, 0x25, 0x0D, 0x0B, 0x03,
	0x5B, 0x08, 0x2B, 0x1B, 0x3B, 0x3A, 0x24, 0x0A, 0x36, 0x41, 0x3C, 0x24,
	0x09, 0x34, 0x2A, 0x13, 0x2A, 0x5D, 0x19, 0x17, 0x02, 0x04, 0x09, 0x32,
	0x02, 0x01, 0x06, 0x1E, 0x19, 0x0D, 0x02, 0x27, 0x02, 0x30, 0x0C, 0x1E,
	0x7A, 0x18, 0x34, 0x04, 0x5E, 0x38, 0x0B, 0x35, 0x2F, 0x39, 0x12, 0x1D,
	0x23, 0x39, 0x58, 0x0B, 0x2A, 0x34, 0x45, 0x20, 0x05, 0x34, 0x25, 0x2A,
	0x02, 0x3A, 0x1C, 0x57, 0x59, 0x27, 0x11, 0x29, 0x57, 0x1A, 0x2D, 0x38,
	0x01, 0x0C, 0x29, 0x27, 0x77, 0x2B, 0x38, 0x0C, 0x2C, 0x3B, 0x5C, 0x0B,
	0x2A, 0x59, 0x34, 0x03, 0x15, 0x05, 0x05, 0x7A, 0x1F, 0x04, 0x2C, 0x12,
	0x6D, 0x1F, 0x00, 0x57, 0x01, 0x26, 0x5B, 0x05, 0x23, 0x02, 0x04, 0x38,
	0x37, 0x06, 0x06, 0x14, 0x19, 0x54, 0x5B, 0x5F, 0x14, 0x5A, 0x0F, 0x14,
	0x31, 0x05, 0x5A, 0x55, 0x56, 0x2E, 0x26, 0x0A, 0x57, 0x18, 0x3C, 0x16,
	0x0D, 0x4A, 0x1D, 0x08, 0x36, 0x28, 0x57, 0x45, 0x5C, 0x24, 0x1D, 0x0F,
	0x05, 0x0F, 0x27, 0x22, 0x25, 0x06, 0x1D, 0x0B, 0x43, 0x32, 0x28, 0x58,
	0x15, 0x5B, 0x39, 0x22, 0x24, 0x7B, 0x14, 0x4E, 0x5D, 0x1D, 0x2E, 0x1E,
	0x00, 0x1F, 0x3B, 0x70, 0x3B, 0x54, 0x2D, 0x0F, 0x38, 0x2D, 0x3B, 0x5F,
	0x26, 0x16, 0x14, 0x58, 0x58, 0x3E, 0x34, 0x35, 0x58, 0x01, 0x44, 0x0D,
	0x34, 0x19, 0x0B, 0x05, 0x17, 0x0B, 0x2C, 0x08, 0x03, 0x27, 0x38, 0x0C,
	0x0A, 0x5C, 0x6D, 0x5D, 0x05, 0x0B, 0x5A, 0x31, 0x0D, 0x56, 0x1A, 0x1D,
	0x05, 0x43, 0x55, 0x03, 0x3F, 0x1A, 0x35, 0x00, 0x5D, 0x06, 0x38, 0x14,
	0x55, 0x59, 0x5E, 0x26, 0x27, 0x56, 0x0B, 0x52, 0x04, 0x1A, 0x18, 0x5D,
	0x52, 0x37, 0x38, 0x07, 0x45, 0x5E, 0x31, 0x09, 0x0C, 0x14, 0x52, 0x34,
	0x19, 0x03, 0x57, 0x3F, 0x2F, 0x0D, 0x50, 0x5C, 0x1C, 0x0B, 0x58, 0x2B,
	0x38, 0x26, 0x21, 0x16, 0x28, 0x14, 0x38, 0x0F, 0x5A, 0x16, 0x0A, 0x59,
	0x28, 0x5C, 0x18, 0x5D, 0x1E, 0x01, 0x05, 0x3B, 0x3B, 0x5B, 0x23, 0x5E,
	0x2D, 0x0C, 0x0F, 0x16, 0x1A, 0x18, 0x26, 0x1F, 0x07, 0x0E, 0x17, 0x5B,
	0x1C, 0x0C, 0x21, 0x03, 0x0C, 0x11, 0x0C, 0x0F, 0x18, 0x2F, 0x27, 0x0E,
	0x04, 0x59, 0x1D, 0x44, 0x75, 0x47, 0x28, 0x00, 0x3F, 0x71, 0x3D, 0x51,
	0x45, 0x03, 0x2D, 0x0F, 0x15, 0x01, 0x01, 0x2B, 0x2E, 0x35, 0x57, 0x5C,
	0x7B, 0x23, 0x36, 0x1C, 0x31, 0x27, 0x18, 0x1B, 0x1D, 0x5D, 0x7A, 0x08,
	0x2A, 0x59, 0x13, 0x73, 0x04, 0x59, 0x14, 0x3C, 0x2C, 0x5B, 0x1B, 0x14,
	0x59, 0x0E, 0x08, 0x0F, 0x14, 0x0A, 0x13, 0x36, 0x31, 0x1D, 0x5D, 0x75,
	0x43, 0x20, 0x22, 0x21, 0x17, 0x15, 0x36, 0x1B, 0x26, 0x35, 0x19, 0x2E,
	0x1C, 0x18, 0x34, 0x55, 0x28, 0x41, 0x3F, 0x23, 0x04, 0x56, 0x34, 0x31,
	0x08, 0x08, 0x32, 0x38, 0x1F, 0x76, 0x1A, 0x32, 0x00, 0x1B, 0x7B, 0x1A,
	0x37, 0x3A, 0x3F, 0x1B, 0x1B, 0x53, 0x0B, 0x59, 0x15, 0x09, 0x54, 0x0C,
	0x26, 0x33, 0x1A, 0x15, 0x06, 0x05, 0x74, 0x3A, 0x50, 0x5A, 0x25, 0x70,
	0x1A, 0x51, 0x1F, 0x53, 0x76, 0x28, 0x11, 0x5C, 0x0A, 0x0A, 0x55, 0x18,
	0x0B, 0x04, 0x23, 0x0A, 0x05, 0x0A, 0x26, 0x77, 0x43, 0x0E, 0x0D, 0x58,
	0x71, 0x34, 0x09, 0x29, 0x00, 0x33, 0x5E, 0x31, 0x3B, 0x19, 0x2D, 0x28,
	0x14, 0x5F, 0x3E, 0x70, 0x19, 0x29, 0x26, 0x5E, 0x0E, 0x5A, 0x15, 0x0B,
	0x32, 0x15, 0x38, 0x22, 0x20, 0x05, 0x1A, 0x1D, 0x59, 0x18, 0x58, 0x28,
	0x0A, 0x38, 0x1E, 0x53, 0x74, 0x43, 0x14, 0x57, 0x1E, 0x05, 0x06, 0x34,
	0x3D, 0x0D, 0x2A, 0x1C, 0x24, 0x2A, 0x05, 0x77, 0x03, 0x12, 0x29, 0x23,
	0x2D, 0x3D, 0x3B, 0x3E, 0x3B, 0x10, 0x1E, 0x14, 0x2A, 0x1F, 0x30, 0x08,
	0x0E, 0x1B, 0x53, 0x36, 0x3F, 0x13, 0x20, 0x22, 0x75, 0x5D, 0x31, 0x59,
	0x1A, 0x3B, 0x2B, 0x25, 0x23, 0x1A, 0x0D, 0x1A, 0x1B, 0x04, 0x33, 0x3A,
	0x21, 0x00, 0x26, 0x24, 0x2A, 0x5F, 0x32, 0x08, 0x26, 0x71, 0x02, 0x55,
	0x3A, 0x09, 0x12, 0x3C, 0x38, 0x59, 0x5A, 0x34, 0x09, 0x37, 0x5D, 0x22,
	0x0B, 0x0B, 0x37, 0x03, 0x5B, 0x16, 0x1F, 0x18, 0x5C, 0x1F, 0x2E, 0x5D,
	0x15, 0x1F, 0x27, 0x72, 0x38, 0x0D, 0x16, 0x1B, 0x7A, 0x35, 0x26, 0x1F,
	0x25, 0x38, 0x35, 0x16, 0x0D, 0x1F, 0x18, 0x19, 0x08, 0x5E, 0x44, 0x12,
	0x29, 0x18, 0x5B, 0x0D, 0x34, 0x23, 0x52, 0x36, 0x05, 0x36, 0x26, 0x50,
	0x39, 0x3B, 0x70, 0x1B, 0x52, 0x1C, 0x1C, 0x08, 0x3E, 0x18, 0x1F, 0x2D,
	0x35, 0x5E, 0x57, 0x21, 0x5B, 0x18, 0x59, 0x2C, 0x0A, 0x01, 0x34, 0x35,
	0x31, 0x22, 0x01, 0x0A, 0x3B, 0x14, 0x1C, 0x53, 0x15, 0x1B, 0x2E, 0x0C,
	0x01, 0x23, 0x09, 0x02, 0x20, 0x3E, 0x2E, 0x1E, 0x58, 0x36, 0x05, 0x20,
	0x35, 0x0E, 0x37, 0x1F, 0x27, 0x14, 0x2D, 0x56, 0x18, 0x0F, 0x24, 0x36,
	0x5A, 0x32, 0x26, 0x5A, 0x34, 0x21, 0x2C, 0x0D, 0x0D, 0x58, 0x1A, 0x1D,
	0x0D, 0x5B, 0x2D, 0x1E, 0x11, 0x76, 0x14, 0x0F, 0x59, 0x03, 0x7B, 0x18,
	0x4E, 0x5F, 0x1B, 0x03, 0x09, 0x0D, 0x1C, 0x1D, 0x27, 0x34, 0x37, 0x01,
	0x53, 0x12, 0x1A, 0x1B, 0x59, 0x38, 0x1B, 0x02, 0x08, 0x1A, 0x5D, 0x17,
	0x2B, 0x2B, 0x23, 0x19, 0x28, 0x2B, 0x53, 0x0F, 0x0F, 0x0F, 0x5C, 0x2A,
	0x0C, 0x33, 0x0A, 0x20, 0x50, 0x0B, 0x2F, 0x2C, 0x18, 0x08, 0x5D, 0x29,
	0x73, 0x2B, 0x2E, 0x5D, 0x08, 0x05, 0x47, 0x56, 0x5D, 0x2E, 0x35, 0x43,
	0x17, 0x14, 0x24, 0x30, 0x14, 0x03, 0x20, 0x11, 0x01, 0x1F, 0x0D, 0x0A,
	0x28, 0x20, 0x0A, 0x37, 0x45, 0x5C, 0x2A, 0x43, 0x17, 0x00, 0x39, 0x32,
	0x3F, 0x2E, 0x41, 0x0E, 0x2A, 0x09, 0x0A, 0x56, 0x18, 0x33, 0x5E, 0x13,
	0x41, 0x0E, 0x14, 0x5F, 0x32, 0x41, 0x1E, 0x04, 0x38, 0x36, 0x5A, 0x3C,
	0x36, 0x28, 0x36, 0x57, 0x31, 0x16, 0x14, 0x0D, 0x5B, 0x06, 0x03, 0x5D,
	0x03, 0x23, 0x28, 0x2F, 0x28, 0x03, 0x0B, 0x38, 0x11, 0x5D, 0x00, 0x5D,
	0x40, 0x6D, 0x2E, 0x06, 0x2C, 0x11, 0x2C, 0x5E, 0x16, 0x5D, 0x3B, 0x30,
	0x06, 0x35, 0x21, 0x06, 0x2F, 0x39, 0x19, 0x57, 0x40, 0x6D, 0x38, 0x0D,
	0x01, 0x3A, 0x29, 0x5E, 0x54, 0x21, 0x20, 0x7B, 0x28, 0x34, 0x0F, 0x32,
	0x20, 0x00, 0x16, 0x41, 0x44, 0x26, 0x35, 0x2E, 0x04, 0x52, 0x0A, 0x20,
	0x2F, 0x3B, 0x0F, 0x11, 0x25, 0x53, 0x20, 0x1D, 0x0A, 0x1E, 0x15, 0x0C,
	0x2C, 0x28, 0x5B, 0x24, 0x5B, 0x28, 0x25, 0x00, 0x52, 0x1C, 0x27, 0x31,
	0x23, 0x29, 0x02, 0x02, 0x15, 0x15, 0x4E, 0x00, 0x08, 0x23, 0x08, 0x17,
	0x3A, 0x11, 0x26, 0x23, 0x32, 0x00, 0x11, 0x23, 0x55, 0x10, 0x2B, 0x11,
	0x74, 0x0A, 0x03, 0x58, 0x5E, 0x2D, 0x0A, 0x24, 0x1B, 0x44, 0x23, 0x22,
	0x0F, 0x1F, 0x53, 0x30, 0x22, 0x29, 0x3D, 0x33, 0x38, 0x27, 0x28, 0x58,
	0x1D, 0x15, 0x1F, 0x12, 0x0B, 0x01, 0x2C, 0x5E, 0x17, 0x3B, 0x0E, 0x30,
	0x54, 0x23, 0x08, 0x5E, 0x2C, 0x39, 0x10, 0x18, 0x00, 0x1B, 0x0A, 0x00,
	0x29, 0x1D, 0x36, 0x24, 0x0F, 0x29, 0x05, 0x2C, 0x5E, 0x26, 0x14, 0x0F,
	0x2E, 0x25, 0x0C, 0x26, 0x2D, 0x34, 0x1D, 0x30, 0x28, 0x52, 0x3A, 0x5E,
	0x3B, 0x24, 0x33, 0x27, 0x27, 0x58, 0x1E, 0x58, 0x08, 0x2F, 0x15, 0x14,
	0x39, 0x1A, 0x20, 0x4E, 0x2F, 0x06, 0x32, 0x03, 0x11, 0x56, 0x0C, 0x2D,
	0x22, 0x25, 0x5B, 0x3E, 0x30, 0x3C, 0x56, 0x5F, 0x08, 0x0D, 0x2E, 0x13,
	0x5D, 0x40, 0x26, 0x07, 0x4A, 0x5F, 0x00, 0x12, 0x2D, 0x58, 0x2D, 0x38,
	0x38, 0x23, 0x53, 0x2A, 0x04, 0x32, 0x09, 0x36, 0x3A, 0x5A, 0x7A, 0x09,
	0x33, 0x1A, 0x09, 0x24, 0x5E, 0x13, 0x5D, 0x39, 0x2D, 0x1F, 0x59, 0x3C,
	0x09, 0x70, 0x59, 0x32, 0x56, 0x44, 0x34, 0x5A, 0x0F, 0x1A, 0x5A, 0x0E,
	0x19, 0x39, 0x5A, 0x53, 0x1B, 0x09, 0x30, 0x3A, 0x25, 0x20, 0x16, 0x07,
	0x58, 0x26, 0x16, 0x5A, 0x05, 0x5B, 0x25, 0x75, 0x43, 0x08, 0x2D, 0x21,
	0x38, 0x5D, 0x52, 0x5F, 0x53, 0x77, 0x1E, 0x2E, 0x5D, 0x0D, 0x06, 0x06,
	0x09, 0x0F, 0x1D, 0x32, 0x5D, 0x2B, 0x45, 0x13, 0x77, 0x23, 0x2D, 0x57,
	0x5A, 0x33, 0x3C, 0x08, 0x3E, 0x04, 0x23, 0x21, 0x0C, 0x0B, 0x44, 0x20,
	0x47, 0x03, 0x2A, 0x39, 0x33, 0x35, 0x17, 0x3B, 0x1D, 0x17, 0x3B, 0x37,
	0x41, 0x22, 0x2F, 0x05, 0x28, 0x18, 0x1E, 0x31, 0x05, 0x56, 0x23, 0x2C,
	0x37, 0x0D, 0x55, 0x5E, 0x1B, 0x0F, 0x35, 0x50, 0x59, 0x25, 0x34, 0x34,
	0x12, 0x3B, 0x05, 0x2D, 0x47, 0x51, 0x04, 0x2F, 0x74, 0x15, 0x58, 0x3E,
	0x09, 0x72, 0x5C, 0x0F, 0x41, 0x1C, 0x2D, 0x55, 0x04, 0x26, 0x29, 0x33,
	0x1A, 0x58, 0x5C, 0x5C, 0x0A, 0x36, 0x11, 0x45, 0x5D, 0x36, 0x39, 0x0E,
	0x59, 0x2F, 0x2C, 0x3A, 0x18, 0x17, 0x0C, 0x3A, 0x39, 0x03, 0x18, 0x39,
	0x21, 0x0E, 0x15, 0x5C, 0x3B, 0x2C, 0x21, 0x14, 0x29, 0x3A, 0x73, 0x1E,
	0x33, 0x36, 0x3C, 0x16, 0x5B, 0x15, 0x1C, 0x07, 0x34, 0x28, 0x00, 0x5B,
	0x11, 0x69, 0x58, 0x14, 0x20, 0x5F, 0x33, 0x07, 0x33, 0x56, 0x0A, 0x10,
	0x43, 0x2B, 0x17, 0x1D, 0x36, 0x18, 0x26, 0x18, 0x1B, 0x2C, 0x04, 0x4E,
	0x45, 0x11, 0x0B, 0x15, 0x05, 0x27, 0x2A, 0x16, 0x3F, 0x35, 0x5B, 0x18,
	0x1B, 0x19, 0x50, 0x36, 0x5E, 0x2C, 0x09, 0x13, 0x41, 0x26, 0x2B, 0x04,
	0x52, 0x20, 0x28, 0x77, 0x1C, 0x3B, 0x5C, 0x1B, 0x0A, 0x3D, 0x51, 0x1F,
	0x1F, 0x27, 0x1D, 0x15, 0x26, 0x27, 0x71, 0x09, 0x00, 0x0A, 0x2F, 0x0C,
	0x03, 0x10, 0x25, 0x24, 0x31, 0x54, 0x0A, 0x5B, 0x03, 0x33, 0x3A, 0x54,
	0x5D, 0x32, 0x12, 0x29, 0x13, 0x0C, 0x40, 0x07, 0x5F, 0x2F, 0x45, 0x52,
	0x27, 0x5A, 0x38, 0x45, 0x40, 0x11, 0x1B, 0x56, 0x14, 0x1E, 0x0A, 0x0E,
	0x19, 0x1F, 0x5C, 0x0D, 0x23, 0x36, 0x0C, 0x24, 0x10, 0x5E, 0x00, 0x3E,
	0x5D, 0x17, 0x3A, 0x2F, 0x3E, 0x1F, 0x73, 0x05, 0x30, 0x23, 0x12, 0x0F,
	0x0E, 0x56, 0x00, 0x5E, 0x28, 0x5F, 0x2A, 0x36, 0x2D, 0x34, 0x59, 0x02,
	0x3A, 0x07, 0x75, 0x39, 0x26, 0x0A, 0x24, 0x30, 0x5E, 0x04, 0x1F, 0x32,
	0x2D, 0x01, 0x07, 0x2C, 0x39, 0x1A, 0x58, 0x17, 0x59, 0x2E, 0x71, 0x26,
	0x27, 0x5E, 0x3E, 0x26, 0x21, 0x08, 0x21, 0x5C, 0x08, 0x18, 0x52, 0x5E,
	0x09, 0x04, 0x2A, 0x34, 0x41, 0x40, 0x75, 0x5E, 0x06, 0x0A, 0x3F, 0x27,
	0x3F, 0x04, 0x56, 0x40, 0x0C, 0x38, 0x0A, 0x45, 0x1E, 0x24, 0x2A, 0x06,
	0x18, 0x52, 0x71, 0x34, 0x15, 0x5F, 0x03, 0x34, 0x25, 0x0C, 0x21, 0x3F,
	0x21, 0x5E, 0x19, 0x29, 0x24, 0x09, 0x09, 0x12, 0x2D, 0x40, 0x71, 0x5E,
	0x56, 0x0B, 0x5C, 0x00, 0x3A, 0x0D, 0x0F, 0x00, 0x7A, 0x55, 0x52, 0x20,
	0x2F, 0x13, 0x43, 0x0F, 0x5D, 0x2F, 0x0D, 0x09, 0x29, 0x2C, 0x06, 0x77,
	0x22, 0x22, 0x05, 0x1B, 0x2C, 0x35, 0x0E, 0x5C, 0x3B, 0x18, 0x0B, 0x54,
	0x1F, 0x25, 0x74, 0x5E, 0x26, 0x5D, 0x06, 0x20, 0x24, 0x53, 0x5B, 0x18,
	0x36, 0x0A, 0x02, 0x2F, 0x1E, 0x24, 0x3A, 0x14, 0x19, 0x06, 0x27, 0x16,
	0x28, 0x3F, 0x25, 0x0A, 0x2E, 0x03, 0x3F, 0x25, 0x2C, 0x18, 0x24, 0x1D,
	0x1F, 0x2A, 0x3C, 0x54, 0x1E, 0x5D, 0x12, 0x47, 0x1B, 0x2B, 0x3F, 0x16,
	0x47, 0x02, 0x0A, 0x53, 0x0F, 0x1F, 0x00, 0x36, 0x59, 0x0D, 0x3E, 0x2F,
	0x01, 0x1B, 0x09, 0x1F, 0x18, 0x56, 0x1F, 0x71, 0x5F, 0x33, 0x5C, 0x3C,
	0x2E, 0x55, 0x02, 0x1B, 0x18, 0x16, 0x3E, 0x59, 0x56, 0x1C, 0x15, 0x15,
	0x58, 0x0A, 0x5D, 0x31, 0x55, 0x02, 0x0A, 0x26, 0x28, 0x16, 0x54, 0x56,
	0x40, 0x08, 0x26, 0x52, 0x45, 0x1D, 0x18, 0x5B, 0x2F, 0x59, 0x27, 0x0E,
	0x1F, 0x30, 0x23, 0x40, 0x17, 0x19, 0x15, 0x17, 0x23, 0x14, 0x5E, 0x4E,
	0x23, 0x58, 0x24, 0x1F, 0x16, 0x5B, 0x31, 0x11, 0x34, 0x54, 0x27, 0x5D,
	0x0D, 0x09, 0x04, 0x5E, 0x1A, 0x37, 0x05, 0x00, 0x1B, 0x1A, 0x08, 0x24,
	0x55, 0x2F, 0x2C, 0x28, 0x2E, 0x4A, 0x3A, 0x08, 0x34, 0x09, 0x53, 0x21,
	0x33, 0x10, 0x5F, 0x52, 0x5E, 0x2C, 0x74, 0x0D, 0x10, 0x36, 0x5B, 0x77,
	0x0F, 0x37, 0x5F, 0x2A, 0x34, 0x06, 0x19, 0x39, 0x07, 0x06, 0x55, 0x35,
	0x0C, 0x31, 0x14, 0x43, 0x19, 0x0F, 0x0F, 0x2F, 0x5C, 0x54, 0x08, 0x26,
	0x70, 0x07, 0x2B, 0x34, 0x0A, 0x0E, 0x59, 0x10, 0x05, 0x3E, 0x7A, 0x26,
	0x14, 0x03, 0x0D, 0x20, 0x22, 0x27, 0x5B, 0x5A, 0x75, 0x55, 0x0E, 0x26,
	0x18, 0x34, 0x0F, 0x18, 0x07, 0x11, 0x07, 0x18, 0x2E, 0x1F, 0x0D, 0x12,
	0x06, 0x53, 0x1B, 0x52, 0x75, 0x1F, 0x0C, 0x5A, 0x03, 0x2B, 0x20, 0x18,
	0x56, 0x3A, 0x7A, 0x18, 0x59, 0x37, 0x05, 0x08, 0x16, 0x57, 0x0C, 0x1A,
	0x23, 0x27, 0x54, 0x5D, 0x3C, 0x3A, 0x1C, 0x57, 0x05, 0x1D, 0x32, 0x28,
	0x56, 0x22, 0x1C, 0x7B, 0x36, 0x07, 0x03, 0x19, 0x14, 0x27, 0x53, 0x05,
	0x20, 0x13, 0x00, 0x4A, 0x3C, 0x1F, 0x30, 0x39, 0x55, 0x2F, 0x07, 0x24,
	0x3C, 0x4A, 0x5F, 0x19, 0x23, 0x1A, 0x0C, 0x5C, 0x38, 0x74, 0x18, 0x2D,
	0x08, 0x5D, 0x13, 0x3B, 0x2B, 0x24, 0x24, 0x27, 0x16, 0x10, 0x27, 0x31,
	0x0A, 0x3B, 0x3B, 0x0A, 0x5C, 0x34, 0x5F, 0x09, 0x00, 0x2D, 0x2F, 0x3C,
	0x2C, 0x0F, 0x1D, 0x34, 0x39, 0x0E, 0x59, 0x23, 0x0A, 0x0B, 0x19, 0x5B,
	0x5E, 0x69, 0x27, 0x11, 0x08, 0x5A, 0x25, 0x5A, 0x58, 0x1D, 0x0E, 0x01,
	0x5B, 0x00, 0x34, 0x3E, 0x77, 0x25, 0x39, 0x1A, 0x5C, 0x7B, 0x1E, 0x26,
	0x21, 0x5E, 0x23, 0x34, 0x29, 0x38, 0x13, 0x72, 0x1F, 0x0C, 0x22, 0x59,
	0x11, 0x3C, 0x2B, 0x00, 0x28, 0x72, 0x1F, 0x1B, 0x57, 0x44, 0x09, 0x1C,
	0x03, 0x5B, 0x1F, 0x33, 0x28, 0x2D, 0x17, 0x52, 0x23, 0x21, 0x28, 0x36,
	0x5D, 0x33, 0x0A, 0x07, 0x1D, 0x59, 0x3A, 0x15, 0x07, 0x0C, 0x0E, 0x70,
	0x2B, 0x59, 0x59, 0x0F, 0x24, 0x16, 0x22, 0x07, 0x11, 0x08, 0x35, 0x57,
	0x5F, 0x3C, 0x72, 0x3C, 0x28, 0x02, 0x1E, 0x24, 0x09, 0x23, 0x26, 0x03,
	0x69, 0x02, 0x35, 0x59, 0x1F, 0x74, 0x18, 0x35, 0x17, 0x3D, 0x14, 0x54,
	0x4E, 0x07, 0x21, 0x01, 0x5C, 0x29, 0x38, 0x0D, 0x3A, 0x3B, 0x0C, 0x14,
	0x24, 0x24, 0x1B, 0x33, 0x5C, 0x1E, 0x11, 0x15, 0x11, 0x09, 0x2E, 0x77,
	0x36, 0x31, 0x0F, 0x05, 0x76, 0x58, 0x15, 0x29, 0x27, 0x2F, 0x01, 0x19,
	0x34, 0x0A, 0x03, 0x0E, 0x58, 0x0C, 0x28, 0x76, 0x19, 0x51, 0x1B, 0x05,
	0x28, 0x06, 0x3B, 0x0A, 0x5C, 0x7A, 0x5A, 0x56, 0x20, 0x44, 0x30, 0x28,
	0x57, 0x23, 0x33, 0x29, 0x06, 0x0E, 0x09, 0x24, 0x23, 0x22, 0x00, 0x2C,
	0x1D, 0x1A, 0x21, 0x25, 0x58, 0x59, 0x7B, 0x0E, 0x51, 0x3E, 0x5E, 0x2C,
	0x3D, 0x58, 0x24, 0x12, 0x34, 0x47, 0x0F, 0x1E, 0x27, 0x1A, 0x43, 0x3B,
	0x3A, 0x0E, 0x75, 0x3A, 0x17, 0x26, 0x21, 0x74, 0x0A, 0x39, 0x2B, 0x32,
	0x0C, 0x34, 0x29, 0x3C, 0x38, 0x08, 0x5E, 0x31, 0x18, 0x0D, 0x32, 0x03,
	0x13, 0x1B, 0x01, 0x73, 0x55, 0x0E, 0x1C, 0x40, 0x2A, 0x20, 0x39, 0x05,
	0x1E, 0x27, 0x25, 0x38, 0x22, 0x0E, 0x36, 0x39, 0x56, 0x58, 0x3F, 0x03,
	0x3F, 0x4A, 0x57, 0x1D, 0x74, 0x59, 0x00, 0x34, 0x00, 0x73, 0x1F, 0x00,
	0x0A, 0x5C, 0x2F, 0x5E, 0x03, 0x18, 0x39, 0x33, 0x58, 0x59, 0x0C, 0x06,
	0x1B, 0x34, 0x27, 0x34, 0x2F, 0x35, 0x08, 0x33, 0x21, 0x0E, 0x36, 0x1F,
	0x07, 0x25, 0x32, 0x31, 0x5E, 0x26, 0x58, 0x1C, 0x20, 0x19, 0x18, 0x1A,
	0x58, 0x30, 0x02, 0x31, 0x0A, 0x1B, 0x12, 0x34, 0x16, 0x02, 0x5F, 0x2C,
	0x08, 0x37, 0x5E, 0x1D, 0x37, 0x1E, 0x0E, 0x00, 0x58, 0x37, 0x38, 0x57,
	0x03, 0x07, 0x26, 0x5E, 0x3B, 0x3E, 0x44, 0x1A, 0x0B, 0x02, 0x39, 0x0D,
	0x75, 0x03, 0x0B, 0x08, 0x0D, 0x73, 0x00, 0x05, 0x21, 0x1E, 0x34, 0x2B,
	0x06, 0x14, 0x2D, 0x17, 0x3F, 0x05, 0x45, 0x5B, 0x33, 0x36, 0x26, 0x2C,
	0x27, 0x15, 0x0E, 0x2F, 0x59, 0x33, 0x70, 0x5A, 0x55, 0x20, 0x5C, 0x70,
	0x39, 0x4A, 0x3C, 0x5B, 0x0A, 0x15, 0x17, 0x1A, 0x1B, 0x33, 0x18, 0x29,
	0x36, 0x12, 0x31, 0x1D, 0x51, 0x2C, 0x2E, 0x69, 0x29, 0x39, 0x3B, 0x05,
	0x05, 0x5C, 0x11, 0x0A, 0x28, 0x36, 0x18, 0x10, 0x0A, 0x0D, 0x2A, 0x35,
	0x0D, 0x24, 0x09, 0x18, 0x1B, 0x08, 0x5F, 0x1E, 0x0E, 0x02, 0x36, 0x1C,
	0x3B, 0x71, 0x1D, 0x19, 0x1F, 0x5B, 0x31, 0x0E, 0x57, 0x5F, 0x08, 0x38,
	0x3E, 0x22, 0x37, 0x21, 0x38, 0x5E, 0x57, 0x3D, 0x0D, 0x30, 0x5D, 0x30,
	0x0F, 0x11, 0x34, 0x0E, 0x54, 0x5D, 0x18, 0x31, 0x09, 0x0B, 0x34, 0x31,
	0x34, 0x55, 0x31, 0x0D, 0x01, 0x38, 0x3D, 0x10, 0x58, 0x05, 0x2A, 0x04,
	0x38, 0x58, 0x3B, 0x73, 0x19, 0x00, 0x05, 0x05, 0x18, 0x14, 0x30, 0x08,
	0x2C, 0x0E, 0x3F, 0x36, 0x1B, 0x03, 0x75, 0x3F, 0x58, 0x05, 0x0A, 0x20,
	0x47, 0x10, 0x5C, 0x27, 0x6D, 0x00, 0x54, 0x3C, 0x1D, 0x2F, 0x43, 0x19,
	0x1E, 0x2D, 0x24, 0x07, 0x39, 0x08, 0x0E, 0x13, 0x09, 0x18, 0x5E, 0x27,
	0x2C, 0x58, 0x30, 0x1D, 0x0D, 0x0D, 0x14, 0x0D, 0x5D, 0x53, 0x2B, 0x59,
	0x25, 0x14, 0x06, 0x2D, 0x15, 0x55, 0x1B, 0x07, 0x32, 0x5A, 0x54, 0x03,
	0x06, 0x00, 0x5E, 0x0E, 0x1E, 0x44, 0x36, 0x5C, 0x59, 0x01, 0x0D, 0x7B,
	0x5D, 0x2A, 0x3D, 0x01, 0x27, 0x5C, 0x50, 0x5E, 0x39, 0x31, 0x14, 0x57,
	0x5B, 0x25, 0x03, 0x06, 0x58, 0x0F, 0x33, 0x2F, 0x0E, 0x28, 0x24, 0x12,
	0x75, 0x1A, 0x2D, 0x2A, 0x1A, 0x74, 0x19, 0x05, 0x58, 0x53, 0x74, 0x0F,
	0x29, 0x16, 0x2E, 0x10, 0x2B, 0x0E, 0x36, 0x13, 0x18, 0x24, 0x4A, 0x1C,
	0x5C, 0x73, 0x0F, 0x26, 0x03, 0x05, 0x10, 0x5A, 0x29, 0x14, 0x29, 0x6D,
	0x43, 0x58, 0x18, 0x27, 0x27, 0x00, 0x04, 0x1E, 0x3E, 0x21, 0x20, 0x54,
	0x39, 0x3A, 0x69, 0x15, 0x53, 0x06, 0x5A, 0x23, 0x3A, 0x07, 0x41, 0x26,
	0x16, 0x29, 0x4A, 0x0A, 0x29, 0x2E, 0x3F, 0x29, 0x20, 0x0D, 0x14, 0x18,
	0x04, 0x57, 0x1E, 0x05, 0x39, 0x15, 0x1B, 0x1D, 0x30, 0x55, 0x2B, 0x0C,
	0x06, 0x28, 0x27, 0x34, 0x5D, 0x20, 0x0E, 0x0A, 0x4A, 0x57, 0x5C, 0x1B,
	0x07, 0x11, 0x0A, 0x27, 0x1A, 0x14, 0x4E, 0x39, 0x1D, 0x12, 0x23, 0x15,
	0x1E, 0x21, 0x0B, 0x5A, 0x10, 0x2D, 0x18, 0x0C, 0x23, 0x0C, 0x3E, 0x5E,
	0x3A, 0x01, 0x4A, 0x41, 0x59, 0x2D, 0x34, 0x12, 0x59, 0x59, 0x7A, 0x18,
	0x10, 0x3D, 0x33, 0x26, 0x28, 0x10, 0x0C, 0x1B, 0x36, 0x1E, 0x33, 0x0F,
	0x1E, 0x23, 0x05, 0x12, 0x2B, 0x3B, 0x70, 0x35, 0x2E, 0x34, 0x23, 0x31,
	0x55, 0x35, 0x5D, 0x03, 0x6D, 0x3F, 0x34, 0x3A, 0x33, 0x30, 0x23, 0x56,
	0x45, 0x09, 0x3A, 0x2A, 0x29, 0x0A, 0x27, 0x14, 0x15, 0x25, 0x38, 0x0D,
	0x01, 0x15, 0x3B, 0x20, 0x0D, 0x2C, 0x0A, 0x10, 0x56, 0x5E, 0x08, 0x3A,
	0x08, 0x14, 0x5F, 0x7A, 0x5B, 0x14, 0x5F, 0x26, 0x2F, 0x0F, 0x52, 0x0C,
	0x0E, 0x21, 0x2A, 0x54, 0x09, 0x26, 0x75, 0x34, 0x04, 0x57, 0x1F, 0x05,
	0x0A, 0x23, 0x22, 0x1A, 0x38, 0x15, 0x34, 0x08, 0x0E, 0x17, 0x3F, 0x15,
	0x21, 0x3F, 0x23, 0x1D, 0x10, 0x57, 0x58, 0x76, 0x1B, 0x52, 0x37, 0x59,
	0x75, 0x19, 0x36, 0x29, 0x1B, 0x04, 0x5B, 0x39, 0x3A, 0x06, 0x75, 0x3F,
	0x03, 0x45, 0x5B, 0x24, 0x02, 0x2F, 0x20, 0x5D, 0x27, 0x23, 0x04, 0x0D,
	0x31, 0x11, 0x2D, 0x0D, 0x07, 0x0D, 0x75, 0x03, 0x0A, 0x2C, 0x26, 0x16,
	0x18, 0x0D, 0x5C, 0x0A, 0x71, 0x21, 0x2D, 0x5E, 0x40, 0x30, 0x22, 0x37,
	0x1E, 0x24, 0x1A, 0x3B, 0x53, 0x3F, 0x3B, 0x11, 0x01, 0x52, 0x02, 0x0A,
	0x36, 0x5F, 0x14, 0x57, 0x18, 0x27, 0x24, 0x28, 0x17, 0x08, 0x71, 0x26,
	0x0D, 0x3D, 0x40, 0x20, 0x0A, 0x53, 0x1A, 0x13, 0x26, 0x20, 0x0F, 0x16,
	0x11, 0x20, 0x2A, 0x31, 0x3F, 0x1E, 0x26, 0x07, 0x33, 0x28, 0x26, 0x01,
	0x2F, 0x56, 0x45, 0x32, 0x16, 0x09, 0x10, 0x03, 0x3A, 0x71, 0x19, 0x05,
	0x5C, 0x0E, 0x14, 0x14, 0x0E, 0x57, 0x5A, 0x15, 0x21, 0x17, 0x45, 0x1B,
	0x73, 0x1C, 0x31, 0x57, 0x01, 0x2A, 0x18, 0x0C, 0x0A, 0x38, 0x71, 0x43,
	0x53, 0x1C, 0x07, 0x29, 0x39, 0x0B, 0x1A, 0x38, 0x29, 0x19, 0x0D, 0x58,
	0x44, 0x27, 0x15, 0x03, 0x04, 0x0E, 0x0C, 0x01, 0x17, 0x5B, 0x58, 0x7B,
	0x19, 0x0E, 0x02, 0x19, 0x08, 0x1A, 0x39, 0x5C, 0x53, 0x09, 0x27, 0x56,
	0x3E, 0x3A, 0x69, 0x54, 0x2E, 0x58, 0x3B, 0x6D, 0x58, 0x39, 0x1C, 0x0D,
	0x76, 0x18, 0x2E, 0x26, 0x12, 0x18, 0x14, 0x1B, 0x27, 0x13, 0x75, 0x43,
	0x05, 0x29, 0x01, 0x1A, 0x21, 0x53, 0x5F, 0x0C, 0x2D, 0x1B, 0x52, 0x59,
	0x19, 0x28, 0x05, 0x32, 0x03, 0x5C, 0x23, 0x27, 0x13, 0x18, 0x58, 0x7A,
	0x5C, 0x52, 0x5D, 0x29, 0x69, 0x23, 0x58, 0x06, 0x0D, 0x30, 0x24, 0x35,
	0x1E, 0x07, 0x0A, 0x55, 0x3B, 0x18, 0x05, 0x75, 0x14, 0x26, 0x02, 0x5B,
	0x30, 0x05, 0x23, 0x41, 0x19, 0x04, 0x5E, 0x19, 0x59, 0x0D, 0x08, 0x00,
	0x51, 0x02, 0x08, 0x33, 0x19, 0x05, 0x2A, 0x09, 0x33, 0x34, 0x50, 0x5C,
	0x1B, 0x77, 0x22, 0x56, 0x3A, 0x2C, 0x21, 0x3C, 0x59, 0x17, 0x3A, 0x38,
	0x09, 0x28, 0x45, 0x0E, 0x28, 0x3F, 0x14, 0x57, 0x1F, 0x16, 0x2E, 0x51,
	0x39, 0x20, 0x77, 0x03, 0x07, 0x20, 0x53, 0x14, 0x5D, 0x2A, 0x14, 0x25,
	0x07, 0x15, 0x05, 0x5D, 0x24, 0x37, 0x5D, 0x39, 0x00, 0x2F, 0x2C, 0x24,
	0x17, 0x3B, 0x06, 0x2B, 0x16, 0x53, 0x20, 0x38, 0x70, 0x1A, 0x4A, 0x0D,
	0x53, 0x3B, 0x15, 0x05, 0x02, 0x0D, 0x36, 0x29, 0x2F, 0x56, 0x0C, 0x75,
	0x1A, 0x26, 0x3F, 0x03, 0x37, 0x38, 0x2F, 0x17, 0x5D, 0x7A, 0x09, 0x19,
	0x3C, 0x0E, 0x27, 0x47, 0x08, 0x5C, 0x59, 0x15, 0x29, 0x0E, 0x1B, 0x27,
	0x26, 0x5D, 0x23, 0x3C, 0x2A, 0x1B, 0x08, 0x24, 0x34, 0x5A, 0x77, 0x09,
	0x0C, 0x57, 0x40, 0x75, 0x18, 0x02, 0x05, 0x31, 0x0A, 0x58, 0x12, 0x18,
	0x5E, 0x0C, 0x0B, 0x13, 0x07, 0x3E, 0x73, 0x3B, 0x33, 0x57, 0x12, 0x7B,
	0x0A, 0x04, 0x5D, 0x21, 0x37, 0x05, 0x29, 0x24, 0x59, 0x74, 0x22, 0x28,
	0x06, 0x5C, 0x7A, 0x22, 0x3B, 0x1F, 0x0A, 0x72, 0x2B, 0x03, 0x3A, 0x1C,
	0x29, 0x21, 0x26, 0x27, 0x04, 0x0E, 0x18, 0x35, 0x14, 0x5A, 0x0E, 0x18,
	0x35, 0x18, 0x33, 0x31, 0x0D, 0x03, 0x26, 0x3F, 0x75, 0x29, 0x56, 0x00,
	0x44, 0x0E, 0x07, 0x58, 0x26, 0x5D, 0x24, 0x1D, 0x34, 0x0B, 0x0A, 0x11,
	0x04, 0x07, 0x37, 0x3F, 0x34, 0x06, 0x35, 0x0A, 0x53, 0x2F, 0x01, 0x22,
	0x16, 0x53, 0x0B, 0x43, 0x4A, 0x05, 0x01, 0x0B, 0x1F, 0x51, 0x5F, 0x06,
	0x12, 0x19, 0x52, 0x17, 0x53, 0x27, 0x3C, 0x1B, 0x58, 0x08, 0x37, 0x38,
	0x13, 0x38, 0x0A, 0x7B, 0x0A, 0x51, 0x07, 0x5E, 0x04, 0x27, 0x4E, 0x0B,
	0x05, 0x16, 0x1A, 0x56, 0x0D, 0x12, 0x34, 0x08, 0x16, 0x20, 0x08, 0x75,
	0x02, 0x56, 0x3C, 0x19, 0x11, 0x3F, 0x52, 0x0D, 0x1F, 0x7B, 0x5E, 0x14,
	0x58, 0x3B, 0x33, 0x34, 0x0E, 0x20, 0x3A, 0x27, 0x5B, 0x55, 0x59, 0x40,
	0x05, 0x38, 0x10, 0x29, 0x3B, 0x12, 0x28, 0x05, 0x01, 0x18, 0x2C, 0x22,
	0x16, 0x16, 0x44, 0x0A, 0x01, 0x2C, 0x19, 0x33, 0x77, 0x1A, 0x05, 0x56,
	0x52, 0x1B, 0x22, 0x00, 0x26, 0x25, 0x37, 0x05, 0x16, 0x36, 0x58, 0x0A,
	0x25, 0x57, 0x0B, 0x53, 0x20, 0x1E, 0x17, 0x1A, 0x40, 0x00, 0x00, 0x09,
	0x3A, 0x59, 0x72, 0x35, 0x56, 0x45, 0x08, 0x69, 0x43, 0x13, 0x3E, 0x0A,
	0x2E, 0x0F, 0x27, 0x04, 0x24, 0x29, 0x39, 0x14, 0x36, 0x2F, 0x69, 0x28,
	0x0F, 0x22, 0x32, 0x29, 0x55, 0x36, 0x17, 0x05, 0x33, 0x29, 0x29, 0x5F,
	0x3C, 0x3B, 0x5F, 0x59, 0x58, 0x25, 0x7B, 0x0B, 0x0F, 0x17, 0x5C, 0x18,
	0x25, 0x29, 0x0B, 0x3F, 0x11, 0x3A, 0x0B, 0x2D, 0x11, 0x24, 0x2A, 0x2D,
	0x34, 0x5C, 0x38, 0x14, 0x07, 0x18, 0x23, 0x0C, 0x07, 0x56, 0x1E, 0x5E,
	0x1B, 0x5C, 0x00, 0x28, 0x29, 0x70, 0x43, 0x0B, 0x2B, 0x19, 0x6D, 0x3A,
	0x4E, 0x3A, 0x39, 0x27, 0x14, 0x18, 0x19, 0x07, 0x10, 0x58, 0x50, 0x0F,
	0x1D, 0x20, 0x01, 0x12, 0x17, 0x09, 0x36, 0x2B, 0x0D, 0x5B, 0x18, 0x71,
	0x39, 0x0F, 0x56, 0x33, 0x18, 0x29, 0x2B, 0x45, 0x44, 0x26, 0x1E, 0x50,
	0x0B, 0x3E, 0x00, 0x0E, 0x52, 0x1A, 0x38, 0x35, 0x58, 0x54, 0x20, 0x3F,
	0x6D, 0x01, 0x0B, 0x3D, 0x07, 0x77, 0x1C, 0x52, 0x41, 0x25, 0x37, 0x09,
	0x37, 0x0C, 0x1E, 0x23, 0x08, 0x31, 0x21, 0x53, 0x33, 0x3C, 0x0F, 0x03,
	0x58, 0x12, 0x2E, 0x08, 0x56, 0x19, 0x20, 0x16, 0x22, 0x08, 0x5E, 0x16,
	0x5E, 0x4A, 0x22, 0x01, 0x24, 0x1B, 0x52, 0x1A, 0x5B, 0x29, 0x43, 0x07,
	0x14, 0x04, 0x0E, 0x54, 0x52, 0x1B, 0x5E, 0x2F, 0x5C, 0x54, 0x1B, 0x25,
	0x10, 0x14, 0x0F, 0x23, 0x06, 0x6D, 0x26, 0x4A, 0x38, 0x18, 0x2C, 0x2B,
	0x27, 0x2D, 0x19, 0x15, 0x43, 0x31, 0x58, 0x22, 0x1A, 0x00, 0x56, 0x14,
	0x0E, 0x74, 0x5B, 0x15, 0x21, 0x18, 0x36, 0x5D, 0x4A, 0x1C, 0x1F, 0x7B,
	0x1C, 0x2E, 0x2C, 0x13, 0x31, 0x14, 0x06, 0x1A, 0x52, 0x23, 0x14, 0x35,
	0x01, 0x08, 0x24, 0x1E, 0x0F, 0x0B, 0x00, 0x69, 0x1B, 0x2B, 0x5A, 0x26,
	0x33, 0x3C, 0x05, 0x38, 0x19, 0x15, 0x28, 0x54, 0x41, 0x0C, 0x32, 0x16,
	0x2F, 0x57, 0x52, 0x75, 0x5C, 0x02, 0x08, 0x2C, 0x17, 0x16, 0x50, 0x39,
	0x11, 0x24, 0x5D, 0x13, 0x5A, 0x1B, 0x20, 0x58, 0x06, 0x26, 0x2D, 0x2C,
	0x07, 0x0E, 0x3E, 0x2C, 0x1A, 0x38, 0x09, 0x22, 0x05, 0x2C, 0x14, 0x32,
	0x5F, 0x23, 0x28, 0x1C, 0x16, 0x34, 0x31, 0x06, 0x2A, 0x14, 0x1A, 0x24,
	0x75, 0x36, 0x0D, 0x19, 0x04, 0x3B, 0x0A, 0x11, 0x1B, 0x08, 0x18, 0x06,
	0x53, 0x1C, 0x11, 0x38, 0x55, 0x0E, 0x41, 0x09, 0x30, 0x16, 0x2C, 0x58,
	0x07, 0x10, 0x47, 0x54, 0x05, 0x2D, 0x33, 0x5A, 0x08, 0x45, 0x19, 0x37,
	0x01, 0x07, 0x26, 0x40, 0x69, 0x0D, 0x12, 0x57, 0x29, 0x26, 0x03, 0x15,
	0x03, 0x52, 0x76, 0x04, 0x2F, 0x5D, 0x5F, 0x2E, 0x35, 0x19, 0x5E, 0x3B,
	0x36, 0x3D, 0x14, 0x5D, 0x05, 0x12, 0x43, 0x02, 0x0B, 0x3E, 0x3A, 0x14,
	0x20, 0x22, 0x07, 0x73, 0x55, 0x13, 0x05, 0x00, 0x2B, 0x5E, 0x32, 0x3E,
	0x02, 0x0D, 0x58, 0x33, 0x5D, 0x0C, 0x0F, 0x34, 0x0B, 0x20, 0x1B, 0x03,
	0x24, 0x03, 0x1E, 0x40, 0x30, 0x3A, 0x39, 0x18, 0x53, 0x0E, 0x27, 0x12,
	0x45, 0x3D, 0x77, 0x26, 0x07, 0x06, 0x3E, 0x2C, 0x5F, 0x11, 0x2A, 0x3E,
	0x34, 0x3E, 0x27, 0x3E, 0x33, 0x0C, 0x0E, 0x0D, 0x5B, 0x52, 0x77, 0x09,
	0x26, 0x1A, 0x32, 0x36, 0x47, 0x50, 0x27, 0x44, 0x0F, 0x01, 0x0C, 0x1E,
	0x1F, 0x21, 0x2A, 0x08, 0x5A, 0x12, 0x04, 0x43, 0x53, 0x18, 0x40, 0x2D,
	0x3C, 0x23, 0x24, 0x05, 0x24, 0x03, 0x35, 0x0F, 0x24, 0x75, 0x1D, 0x18,
	0x5D, 0x2C, 0x24, 0x22, 0x58, 0x29, 0x33, 0x7B, 0x38, 0x11, 0x37, 0x5D,
	0x00, 0x38, 0x58, 0x39, 0x04, 0x70, 0x20, 0x27, 0x1E, 0x39, 0x17, 0x34,
	0x39, 0x1B, 0x0C, 0x7A, 0x1A, 0x29, 0x1B, 0x1B, 0x76, 0x14, 0x04, 0x1E,
	0x08, 0x00, 0x2E, 0x54, 0x18, 0x1E, 0x37, 0x05, 0x4A, 0x24, 0x5B, 0x20,
	0x3C, 0x27, 0x0F, 0x1A, 0x36, 0x0A, 0x13, 0x04, 0x32, 0x07, 0x06, 0x16,
	0x3A, 0x0A, 0x30, 0x1B, 0x36, 0x5A, 0x26, 0x6D, 0x06, 0x17, 0x5B, 0x25,
	0x12, 0x09, 0x0A, 0x0D, 0x25, 0x0A, 0x05, 0x2B, 0x37, 0x3E, 0x18, 0x06,
	0x08, 0x00, 0x0D, 0x01, 0x5C, 0x2A, 0x02, 0x27, 0x1A, 0x23, 0x2A, 0x1B,
	0x3F, 0x69, 0x3B, 0x09, 0x24, 0x0E, 0x2C, 0x18, 0x12, 0x1D, 0x03, 0x04,
	0x3D, 0x56, 0x08, 0x5B, 0x31, 0x09, 0x13, 0x1B, 0x5A, 0x2F, 0x5B, 0x4E,
	0x21, 0x44, 0x0D, 0x01, 0x2E, 0x19, 0x58, 0x24, 0x39, 0x16, 0x5F, 0x05,
	0x0A, 0x43, 0x35, 0x03, 0x13, 0x11, 0x59, 0x4A, 0x07, 0x3F, 0x74, 0x0D,
	0x4A, 0x06, 0x13, 0x0C, 0x0E, 0x51, 0x0D, 0x3D, 0x37, 0x3F, 0x3B, 0x5C,
	0x12, 0x26, 0x59, 0x53, 0x0A, 0x13, 0x69, 0x15, 0x17, 0x1E, 0x0E, 0x72,
	0x1E, 0x31, 0x56, 0x00, 0x0F, 0x1C, 0x30, 0x19, 0x02, 0x69, 0x1C, 0x55,
	0x5C, 0x3B, 0x10, 0x02, 0x39, 0x28, 0x01, 0x13, 0x00, 0x25, 0x2B, 0x07,
	0x05, 0x19, 0x35, 0x1B, 0x13, 0x17, 0x3F, 0x0F, 0x37, 0x20, 0x72, 0x06,
	0x29, 0x36, 0x3F, 0x06, 0x24, 0x16, 0x17, 0x5A, 0x24, 0x55, 0x32, 0x0A,
	0x02, 0x34, 0x29, 0x0D, 0x2A, 0x19, 0x2C, 0x01, 0x0F, 0x39, 0x1D, 0x16,
	0x5B, 0x39, 0x34, 0x11, 0x29, 0x08, 0x39, 0x14, 0x40, 0x27, 0x3D, 0x55,
	0x3A, 0x0A, 0x0B, 0x1F, 0x07, 0x00, 0x3B, 0x00, 0x54, 0x53, 0x56, 0x06,
	0x24, 0x01, 0x2E, 0x2B, 0x19, 0x1B, 0x16, 0x2B, 0x18, 0x5A, 0x1B, 0x38,
	0x53, 0x36, 0x04, 0x36, 0x1E, 0x57, 0x59, 0x3B, 0x71, 0x3B, 0x58, 0x05,
	0x58, 0x6D, 0x26, 0x59, 0x0C, 0x59, 0x30, 0x5C, 0x23, 0x27, 0x0E, 0x0D,
	0x5F, 0x02, 0x0D, 0x26, 0x24, 0x16, 0x52, 0x3B, 0x3A, 0x26, 0x43, 0x2A,
	0x41, 0x58, 0x2D, 0x2E, 0x14, 0x37, 0x29, 0x33, 0x5D, 0x52, 0x45, 0x40,
	0x6D, 0x08, 0x16, 0x5C, 0x04, 0x32, 0x1B, 0x04, 0x19, 0x1B, 0x14, 0x5F,
	0x36, 0x5B, 0x20, 0x15, 0x3F, 0x34, 0x3E, 0x05, 0x10, 0x2B, 0x19, 0x41,
	0x3C, 0x26, 0x5A, 0x09, 0x0F, 0x0E, 0x3B, 0x23, 0x16, 0x37, 0x5E, 0x3A,
	0x3A, 0x29, 0x2D, 0x19, 0x35, 0x5E, 0x56, 0x1C, 0x31, 0x72, 0x0F, 0x2C,
	0x5D, 0x58, 0x69, 0x02, 0x0C, 0x3B, 0x59, 0x1B, 0x55, 0x30, 0x5A, 0x12,
	0x0B, 0x54, 0x08, 0x3C, 0x0D, 0x09, 0x5C, 0x4E, 0x41, 0x24, 0x34, 0x1C,
	0x33, 0x41, 0x08, 0x33, 0x3C, 0x32, 0x1F, 0x1F, 0x3B, 0x36, 0x23, 0x20,
	0x3E, 0x74, 0x02, 0x29, 0x04, 0x33, 0x0F, 0x23, 0x0B, 0x57, 0x38, 0x75,
	0x54, 0x24, 0x07, 0x11, 0x74, 0x3D, 0x08, 0x1F, 0x0A, 0x07, 0x0D, 0x52,
	0x16, 0x2F, 0x69, 0x15, 0x59, 0x06, 0x5A, 0x12, 0x34, 0x22, 0x5B, 0x53,
	0x34, 0x19, 0x1B, 0x21, 0x26, 0x1A, 0x27, 0x52, 0x59, 0x04, 0x29, 0x34,
	0x54, 0x59, 0x5C, 0x72, 0x43, 0x0F, 0x16, 0x13, 0x0E, 0x3B, 0x58, 0x25,
	0x00, 0x72, 0x2E, 0x0F, 0x1D, 0x05, 0x71, 0x3B, 0x51, 0x24, 0x2D, 0x12,
	0x5E, 0x0E, 0x5C, 0x58, 0x70, 0x02, 0x52, 0x59, 0x52, 0x08, 0x1E, 0x52,
	0x27, 0x58, 0x0D, 0x03, 0x12, 0x25, 0x26, 0x06, 0x47, 0x36, 0x0F, 0x1D,
	0x07, 0x02, 0x0B, 0x08, 0x25, 0x33, 0x5C, 0x2A, 0x03, 0x0D, 0x1A, 0x55,
	0x2A, 0x04, 0x07, 0x31, 0x01, 0x02, 0x00, 0x5B, 0x32, 0x18, 0x2F, 0x0B,
	0x25, 0x0D, 0x24, 0x31, 0x28, 0x25, 0x3B, 0x1F, 0x58, 0x56, 0x24, 0x20,
	0x18, 0x31, 0x16, 0x31, 0x27, 0x05, 0x07, 0x26, 0x0A, 0x72, 0x3C, 0x4E,
	0x14, 0x0A, 0x0D, 0x0E, 0x33, 0x18, 0x1D, 0x05, 0x59, 0x27, 0x23, 0x3F,
	0x75, 0x09, 0x31, 0x26, 0x5A, 0x28, 0x18, 0x17, 0x5E, 0x0A, 0x37, 0x43,
	0x53, 0x23, 0x0F, 0x72, 0x47, 0x03, 0x06, 0x05, 0x32, 0x23, 0x31, 0x59,
	0x23, 0x1B, 0x19, 0x14, 0x3D, 0x23, 0x36, 0x5F, 0x2D, 0x36, 0x05, 0x23,
	0x36, 0x36, 0x3C, 0x3F, 0x0F, 0x03, 0x19, 0x56, 0x09, 0x26, 0x0E, 0x17,
	0x05, 0x26, 0x14, 0x20, 0x51, 0x57, 0x06, 0x20, 0x05, 0x4E, 0x1E, 0x23,
	0x36, 0x05, 0x17, 0x0C, 0x3A, 0x7A, 0x5C, 0x38, 0x0B, 0x11, 0x27, 0x14,
	0x58, 0x5F, 0x3F, 0x24, 0x5A, 0x16, 0x0A, 0x59, 0x71, 0x5E, 0x12, 0x3D,
	0x06, 0x34, 0x5A, 0x05, 0x3A, 0x23, 0x12, 0x35, 0x26, 0x07, 0x21, 0x0C,
	0x1A, 0x05, 0x04, 0x1C, 0x30, 0x22, 0x53, 0x5C, 0x29, 0x2A, 0x5B, 0x58,
	0x37, 0x53, 0x2E, 0x18, 0x17, 0x20, 0x28, 0x13, 0x2A, 0x52, 0x58, 0x5C,
	0x1A, 0x18, 0x52, 0x08, 0x2D, 0x00, 0x36, 0x18, 0x5A, 0x08, 0x25, 0x2A,
	0x10, 0x00, 0x5A, 0x16, 0x28, 0x59, 0x3E, 0x33, 0x33, 0x3A, 0x4E, 0x08,
	0x01, 0x0A, 0x55, 0x4E, 0x0F, 0x5F, 0x71, 0x0E, 0x04, 0x3F, 0x3B, 0x33,
	0x3A, 0x38, 0x21, 0x12, 0x33, 0x5A, 0x39, 0x3A, 0x5C, 0x05, 0x35, 0x0C,
	0x26, 0x01, 0x0E, 0x36, 0x17, 0x38, 0x0C, 0x6D, 0x02, 0x33, 0x16, 0x01,
	0x2E, 0x18, 0x53, 0x08, 0x20, 0x0A, 0x5A, 0x16, 0x23, 0x38, 0x12, 0x59,
	0x52, 0x0F, 0x23, 0x18, 0x1A, 0x3B, 0x5B, 0x39, 0x32, 0x59, 0x10, 0x07,
	0x33, 0x25, 0x59, 0x35, 0x24, 0x40, 0x38, 0x43, 0x14, 0x3E, 0x08, 0x06,
	0x36, 0x03, 0x2A, 0x28, 0x2C, 0x2A, 0x13, 0x1E, 0x5B, 0x75, 0x2A, 0x13,
	0x14, 0x0C, 0x30, 0x1D, 0x0B, 0x21, 0x01, 0x0A, 0x1B, 0x2C, 0x5A, 0x52,
	0x16, 0x0F, 0x04, 0x3C, 0x3A, 0x21, 0x07, 0x1B, 0x01, 0x52, 0x0F, 0x0A,
	0x0A, 0x45, 0x3D, 0x28, 0x38, 0x11, 0x01, 0x08, 0x04, 0x01, 0x59, 0x09,
	0x12, 0x06, 0x29, 0x4A, 0x03, 0x44, 0x75, 0x0D, 0x55, 0x0C, 0x20, 0x72,
	0x16, 0x51, 0x22, 0x3B, 0x6D, 0x0F, 0x15, 0x3A, 0x23, 0x71, 0x3F, 0x08,
	0x28, 0x07, 0x75, 0x35, 0x52, 0x41, 0x03, 0x0E, 0x02, 0x2F, 0x45, 0x0F,
	0x7B, 0x35, 0x55, 0x21, 0x0C, 0x1A, 0x5C, 0x0C, 0x14, 0x28, 0x09, 0x24,
	0x52, 0x5A, 0x01, 0x12, 0x1F, 0x0C, 0x5C, 0x1B, 0x12, 0x0A, 0x03, 0x5F,
	0x5C, 0x03, 0x47, 0x13, 0x06, 0x07, 0x12, 0x5A, 0x54, 0x27, 0x08, 0x77,
	0x09, 0x0B, 0x20, 0x23, 0x2C, 0x34, 0x33, 0x0A, 0x1D, 0x0A, 0x34, 0x22,
	0x02, 0x24, 0x1A, 0x18, 0x0D, 0x18, 0x07, 0x11, 0x02, 0x16, 0x16, 0x5B,
	0x7B, 0x24, 0x54, 0x0D, 0x02, 0x36, 0x43, 0x16, 0x1D, 0x0D, 0x0D, 0x00,
	0x11, 0x1B, 0x09, 0x69, 0x15, 0x59, 0x03, 0x01, 0x27, 0x00, 0x10, 0x3D,
	0x23, 0x77, 0x07, 0x56, 0x5D, 0x53, 0x35, 0x47, 0x07, 0x26, 0x25, 0x07,
	0x58, 0x2C, 0x1F, 0x06, 0x32, 0x2B, 0x56, 0x16, 0x3D, 0x24, 0x54, 0x35,
	0x5E, 0x52, 0x76, 0x5F, 0x07, 0x58, 0x32, 0x73, 0x16, 0x56, 0x1C, 0x13,
	0x69, 0x3D, 0x27, 0x3B, 0x1F, 0x74, 0x07, 0x2F, 0x1C, 0x02, 0x3B, 0x34,
	0x29, 0x22, 0x04, 0x6D, 0x27, 0x07, 0x02, 0x3C, 0x70, 0x2B, 0x52, 0x1E,
	0x39, 0x34, 0x20, 0x24, 0x1E, 0x0A, 0x0A, 0x5D, 0x35, 0x08, 0x1E, 0x15,
	0x06, 0x34, 0x57, 0x1E, 0x6D, 0x3B, 0x25, 0x1A, 0x1B, 0x32, 0x1B, 0x53,
	0x1E, 0x2E, 0x0A, 0x35, 0x57, 0x41, 0x2E, 0x06, 0x28, 0x53, 0x5B, 0x0E,
	0x73, 0x00, 0x25, 0x14, 0x5B, 0x37, 0x5F, 0x0C, 0x37, 0x52, 0x0D, 0x03,
	0x0F, 0x03, 0x1D, 0x75, 0x08, 0x0F, 0x59, 0x3A, 0x74, 0x0F, 0x2E, 0x03,
	0x11, 0x12, 0x23, 0x26, 0x03, 0x40, 0x69, 0x06, 0x20, 0x5C, 0x3F, 0x21,
	0x1D, 0x4A, 0x25, 0x29, 0x70, 0x1B, 0x4E, 0x20, 0x0E, 0x28, 0x43, 0x56,
	0x0B, 0x1D, 0x33, 0x2E, 0x59, 0x0F, 0x08, 0x26, 0x15, 0x2B, 0x3B, 0x06,
	0x24, 0x1E, 0x24, 0x39, 0x12, 0x76, 0x22, 0x04, 0x0C, 0x3F, 0x6D, 0x0F,
	0x51, 0x1C, 0x23, 0x0E, 0x04, 0x0B, 0x45, 0x1B, 0x2D, 0x3C, 0x36, 0x36,
	0x05, 0x28, 0x38, 0x07, 0x5E, 0x05, 0x12, 0x0D, 0x54, 0x5E, 0x2D, 0x0C,
	0x1E, 0x29, 0x3E, 0x0D, 0x2C, 0x2F, 0x04, 0x18, 0x5C, 0x31, 0x5C, 0x51,
	0x56, 0x11, 0x34, 0x58, 0x12, 0x5F, 0x1E, 0x17, 0x47, 0x3B, 0x5E, 0x52,
	0x23, 0x43, 0x10, 0x5B, 0x00, 0x14, 0x0E, 0x1B, 0x41, 0x00, 0x77, 0x35,
	0x2E, 0x41, 0x03, 0x17, 0x5B, 0x14, 0x27, 0x12, 0x76, 0x01, 0x14, 0x29,
	0x5D, 0x01, 0x55, 0x10, 0x1E, 0x5A, 0x0A, 0x0F, 0x08, 0x57, 0x2F, 0x08,
	0x27, 0x16, 0x5E, 0x09, 0x1A, 0x35, 0x14, 0x3E, 0x23, 0x37, 0x04, 0x4E,
	0x00, 0x44, 0x3A, 0x5A, 0x03, 0x3B, 0x27, 0x76, 0x1E, 0x04, 0x3C, 0x06,
	0x73, 0x16, 0x19, 0x29, 0x5C, 0x03, 0x1B, 0x51, 0x58, 0x38, 0x76, 0x0B,
	0x3B, 0x56, 0x59, 0x74, 0x2B, 0x31, 0x26, 0x52, 0x75, 0x1C, 0x16, 0x3E,
	0x11, 0x2D, 0x09, 0x15, 0x20, 0x19, 0x75, 0x22, 0x52, 0x3B, 0x11, 0x32,
	0x5A, 0x19, 0x0A, 0x3D, 0x24, 0x28, 0x05, 0x5F, 0x3B, 0x71, 0x16, 0x12,
	0x22, 0x52, 0x74, 0x5B, 0x20, 0x5A, 0x32, 0x24, 0x15, 0x2D, 0x3F, 0x0E,
	0x37, 0x16, 0x07, 0x26, 0x25, 0x2E, 0x03, 0x18, 0x25, 0x23, 0x2C, 0x06,
	0x54, 0x1C, 0x31, 0x2C, 0x5C, 0x16, 0x0B, 0x38, 0x13, 0x3F, 0x02, 0x29,
	0x3B, 0x29, 0x43, 0x04, 0x45, 0x52, 0x2E, 0x1B, 0x16, 0x45, 0x24, 0x08,
	0x2E, 0x06, 0x45, 0x28, 0x16, 0x5D, 0x23, 0x58, 0x07, 0x6D, 0x1B, 0x10,
	0x19, 0x59, 0x0D, 0x06, 0x13, 0x05, 0x3C, 0x7A, 0x0F, 0x2D, 0x19, 0x1A,
	0x21, 0x22, 0x2E, 0x07, 0x1E, 0x2F, 0x08, 0x10, 0x3A, 0x53, 0x7A, 0x0D,
	0x4E, 0x45, 0x02, 0x0D, 0x54, 0x36, 0x1B, 0x39, 0x7B, 0x16, 0x34, 0x07,
	0x06, 0x20, 0x3F, 0x50, 0x23, 0x3B, 0x01, 0x36, 0x10, 0x0F, 0x5E, 0x0A,
	0x2F, 0x34, 0x5E, 0x5C, 0x32, 0x19, 0x34, 0x1D, 0x1E, 0x17, 0x22, 0x3B,
	0x3A, 0x2E, 0x28, 0x38, 0x14, 0x2A, 0x19, 0x2D, 0x0F, 0x0E, 0x22, 0x09,
	0x3B, 0x2D, 0x31, 0x59, 0x53, 0x69, 0x54, 0x50, 0x1E, 0x09, 0x1B, 0x02,
	0x36, 0x1F, 0x00, 0x71, 0x09, 0x26, 0x36, 0x5B, 0x77, 0x47, 0x2B, 0x5B,
	0x02, 0x3A, 0x5E, 0x22, 0x00, 0x5F, 0x35, 0x0B, 0x52, 0x5C, 0x3F, 0x17,
	0x19, 0x4E, 0x3A, 0x53, 0x24, 0x1C, 0x22, 0x1B, 0x0F, 0x15, 0x1A, 0x13,
	0x2B, 0x2E, 0x0A, 0x2B, 0x3B, 0x45, 0x19, 0x7B, 0x14, 0x4A, 0x58, 0x31,
	0x27, 0x1B, 0x39, 0x5B, 0x20, 0x3B, 0x36, 0x17, 0x03, 0x11, 0x35, 0x5C,
	0x4E, 0x0F, 0x26, 0x0C, 0x5D, 0x36, 0x5B, 0x24, 0x00, 0x47, 0x12, 0x21,
	0x5A, 0x71, 0x1C, 0x17, 0x5F, 0x31, 0x3A, 0x55, 0x02, 0x39, 0x29, 0x6D,
	0x5A, 0x57, 0x03, 0x00, 0x69, 0x35, 0x53, 0x45, 0x19, 0x26, 0x58, 0x50,
	0x1B, 0x2F, 0x74, 0x0B, 0x18, 0x41, 0x3C, 0x2A, 0x28, 0x52, 0x19, 0x19,
	0x36, 0x0F, 0x0B, 0x2B, 0x24, 0x1B, 0x0F, 0x26, 0x2D, 0x5A, 0x7A, 0x09,
	0x12, 0x04, 0x18, 0x35, 0x54, 0x29, 0x36, 0x33, 0x2D, 0x08, 0x0C, 0x1B,
	0x07, 0x0C, 0x07, 0x00, 0x1F, 0x1F, 0x15, 0x0D, 0x07, 0x39, 0x3D, 0x6D,
	0x29, 0x53, 0x3E, 0x0A, 0x3A, 0x20, 0x30, 0x41, 0x1D, 0x1B, 0x04, 0x12,
	0x29, 0x1B, 0x0B, 0x58, 0x03, 0x1A, 0x0D, 0x08, 0x55, 0x28, 0x3B, 0x24,
	0x12, 0x15, 0x04, 0x21, 0x0E, 0x3B, 0x3A, 0x11, 0x3D, 0x27, 0x20, 0x06,
	0x14, 0x3F, 0x5A, 0x33, 0x00, 0x4E, 0x39, 0x53, 0x71, 0x59, 0x59, 0x00,
	0x1E, 0x38, 0x01, 0x2E, 0x29, 0x39, 0x36, 0x27, 0x17, 0x08, 0x21, 0x24,
	0x43, 0x2F, 0x27, 0x18, 0x36, 0x55, 0x34, 0x57, 0x52, 0x21, 0x1F, 0x19,
	0x01, 0x1B, 0x69, 0x02, 0x08, 0x56, 0x0C, 0x69, 0x23, 0x13, 0x5A, 0x3C,
	0x32, 0x03, 0x03, 0x0C, 0x1F, 0x33, 0x03, 0x2F, 0x0B, 0x44, 0x08, 0x2D,
	0x52, 0x23, 0x24, 0x21, 0x0E, 0x27, 0x3E, 0x00, 0x27, 0x01, 0x0F, 0x39,
	0x1C, 0x38, 0x5F, 0x0C, 0x17, 0x44, 0x37, 0x58, 0x39, 0x3B, 0x5C, 0x7B,
	0x02, 0x0A, 0x04, 0x1F, 0x0C, 0x28, 0x15, 0x14, 0x18, 0x69, 0x2E, 0x3B,
	0x14, 0x25, 0x23, 0x2D, 0x2E, 0x5A, 0x38, 0x2C, 0x36, 0x38, 0x08, 0x0F,
	0x18, 0x23, 0x57, 0x39, 0x22, 0x10, 0x19, 0x07, 0x03, 0x5F, 0x6D, 0x43,
	0x10, 0x2A, 0x24, 0x15, 0x39, 0x2B, 0x18, 0x32, 0x73, 0x58, 0x55, 0x3B,
	0x44, 0x2A, 0x07, 0x51, 0x14, 0x05, 0x34, 0x1C, 0x34, 0x01, 0x1E, 0x73,
	0x14, 0x2B, 0x27, 0x1E, 0x1A, 0x38, 0x4A, 0x21, 0x1B, 0x36, 0x0D, 0x02,
	0x3A, 0x5A, 0x37, 0x54, 0x03, 0x22, 0x39, 0x08, 0x05, 0x1B, 0x5D, 0x13,
	0x28, 0x3B, 0x18, 0x41, 0x0D, 0x16, 0x1C, 0x2B, 0x03, 0x19, 0x29, 0x08,
	0x14, 0x22, 0x1D, 0x32, 0x1C, 0x2B, 0x0A, 0x0D, 0x38, 0x21, 0x54, 0x0C,
	0x19, 0x24, 0x00, 0x29, 0x1B, 0x5E, 0x0A, 0x29, 0x39, 0x57, 0x3F, 0x11,
	0x2F, 0x03, 0x0A, 0x5A, 0x74, 0x1C, 0x4E, 0x18, 0x2D, 0x75, 0x1A, 0x59,
	0x5A, 0x31, 0x00, 0x0F, 0x00, 0x1A, 0x2C, 0x2D, 0x26, 0x33, 0x1B, 0x1B,
	0x2A, 0x5D, 0x53, 0x18, 0x38, 0x71, 0x5C, 0x27, 0x39, 0x5E, 0x74, 0x5D,
	0x14, 0x3B, 0x06, 0x0D, 0x06, 0x22, 0x5F, 0x1B, 0x72, 0x43, 0x0C, 0x34,
	0x58, 0x21, 0x0B, 0x23, 0x28, 0x5D, 0x69, 0x5E, 0x25, 0x08, 0x1E, 0x28,
	0x2A, 0x53, 0x03, 0x1F, 0x69, 0x3B, 0x09, 0x5F, 0x59, 0x0E, 0x2D, 0x0C,
	0x20, 0x05, 0x23, 0x5B, 0x3B, 0x1A, 0x5D, 0x1B, 0x20, 0x22, 0x03, 0x02,
	0x7B, 0x1D, 0x0E, 0x41, 0x58, 0x75, 0x5B, 0x53, 0x17, 0x3B, 0x03, 0x1C,
	0x03, 0x5D, 0x27, 0x73, 0x09, 0x10, 0x39, 0x3E, 0x34, 0x05, 0x33, 0x04,
	0x11, 0x69, 0x5E, 0x19, 0x2A, 0x07, 0x0D, 0x5F, 0x14, 0x14, 0x3F, 0x28,
	0x59, 0x14, 0x39, 0x27, 0x30, 0x14, 0x05, 0x29, 0x00, 0x0A, 0x01, 0x31,
	0x18, 0x5D, 0x35, 0x3C, 0x14, 0x5D, 0x3F, 0x24, 0x0E, 0x29, 0x3A, 0x5B,
	0x74, 0x5D, 0x50, 0x2C, 0x23, 0x72, 0x1D, 0x11, 0x09, 0x29, 0x26, 0x0A,
	0x16, 0x14, 0x5B, 0x7B, 0x02, 0x0B, 0x58, 0x20, 0x24, 0x38, 0x19, 0x57,
	0x19, 0x36, 0x59, 0x09, 0x3C, 0x24, 0x2F, 0x54, 0x15, 0x04, 0x26, 0x69,
	0x00, 0x56, 0x04, 0x5C, 0x69, 0x34, 0x09, 0x06, 0x2F, 0x3B, 0x21, 0x05,
	0x1A, 0x33, 0x2B, 0x15, 0x00, 0x29, 0x12, 0x16, 0x05, 0x38, 0x28, 0x19,
	0x12, 0x1D, 0x50, 0x3E, 0x28, 0x34, 0x58, 0x4A, 0x0A, 0x1A, 0x2A, 0x2B,
	0x2E, 0x3A, 0x33, 0x08, 0x58, 0x34, 0x5B, 0x31, 0x28, 0x14, 0x22, 0x0C,
	0x1A, 0x18, 0x3B, 0x14, 0x1D, 0x3C, 0x21, 0x2B, 0x2E, 0x06, 0x07, 0x16,
	0x2A, 0x1B, 0x5B, 0x00, 0x73, 0x43, 0x15, 0x5B, 0x32, 0x69, 0x54, 0x0D,
	0x17, 0x53, 0x1A, 0x0E, 0x04, 0x03, 0x1C, 0x74, 0x07, 0x0A, 0x2B, 0x40,
	0x2F, 0x5C, 0x2A, 0x23, 0x44, 0x0A, 0x24, 0x34, 0x0C, 0x1D, 0x09, 0x1D,
	0x06, 0x0B, 0x2C, 0x3A, 0x0B, 0x0D, 0x39, 0x1D, 0x33, 0x21, 0x0C, 0x36,
	0x2D, 0x2A, 0x5F, 0x4E, 0x1D, 0x3C, 0x3B, 0x0D, 0x02, 0x41, 0x25, 0x0C,
	0x55, 0x3B, 0x18, 0x33, 0x23, 0x5E, 0x54, 0x24, 0x0F, 0x16, 0x34, 0x00,
	0x01, 0x3B, 0x2E, 0x16, 0x0B, 0x21, 0x3F, 0x1B, 0x1D, 0x23, 0x03, 0x2D,
	0x2D, 0x5F, 0x35, 0x1B, 0x3F, 0x3B, 0x28, 0x15, 0x1E, 0x2C, 0x6D, 0x23,
	0x2D, 0x5F, 0x01, 0x76, 0x18, 0x12, 0x1B, 0x3B, 0x0B, 0x0E, 0x16, 0x08,
	0x12, 0x77, 0x55, 0x30, 0x1E, 0x29, 0x7B, 0x1A, 0x4A, 0x5A, 0x39, 0x71,
	0x3A, 0x12, 0x57, 0x05, 0x3A, 0x01, 0x19, 0x2A, 0x58, 0x7A, 0x55, 0x0C,
	0x0A, 0x20, 0x04, 0x3B, 0x31, 0x3E, 0x11, 0x17, 0x09, 0x02, 0x2D, 0x1E,
	0x3B, 0x3A, 0x07, 0x26, 0x1F, 0x14, 0x43, 0x51, 0x18, 0x0E, 0x24, 0x2D,
	0x39, 0x22, 0x21, 0x18, 0x54, 0x2B, 0x08, 0x59, 0x7B, 0x5A, 0x2E, 0x39,
	0x0E, 0x77, 0x22, 0x09, 0x27, 0x59, 0x0E, 0x06, 0x4E, 0x2F, 0x11, 0x08,
	0x16, 0x59, 0x5D, 0x0A, 0x05, 0x3F, 0x02, 0x00, 0x0F, 0x36, 0x25, 0x03,
	0x28, 0x23, 0x1B, 0x58, 0x35, 0x45, 0x22, 0x18, 0x3D, 0x2F, 0x05, 0x5B,
	0x2C, 0x19, 0x30, 0x39, 0x23, 0x2C, 0x26, 0x28, 0x0B, 0x52, 0x0E, 0x0D,
	0x30, 0x3F, 0x23, 0x16, 0x24, 0x37, 0x0B, 0x39, 0x17, 0x47, 0x17, 0x00,
	0x27, 0x23, 0x59, 0x4E, 0x23, 0x58, 0x04, 0x59, 0x0D, 0x56, 0x06, 0x16,
	0x1E, 0x0F, 0x3A, 0x44, 0x71, 0x25, 0x19, 0x0D, 0x59, 0x3A, 0x14, 0x58,
	0x28, 0x05, 0x3A, 0x5D, 0x28, 0x57, 0x1F, 0x2F, 0x34, 0x28, 0x1D, 0x5F,
	0x12, 0x05, 0x2E, 0x25, 0x59, 0x36, 0x21, 0x38, 0x5B, 0x0F, 0x1B, 0x5B,
	0x0F, 0x1C, 0x2F, 0x76, 0x3E, 0x02, 0x58, 0x22, 0x7B, 0x0F, 0x54, 0x1E,
	0x3C, 0x7A, 0x04, 0x54, 0x58, 0x13, 0x23, 0x19, 0x14, 0x34, 0x27, 0x0A,
	0x54, 0x52, 0x5C, 0x0F, 0x6D, 0x01, 0x52, 0x18, 0x5A, 0x71, 0x08, 0x15,
	0x17, 0x33, 0x06, 0x1A, 0x4E, 0x09, 0x31, 0x7B, 0x2F, 0x22, 0x22, 0x01,
	0x21, 0x0F, 0x14, 0x04, 0x58, 0x35, 0x5A, 0x29, 0x2A, 0x20, 0x14, 0x19,
	0x10, 0x5A, 0x44, 0x33, 0x5A, 0x04, 0x5E, 0x3A, 0x71, 0x47, 0x56, 0x28,
	0x06, 0x12, 0x21, 0x19, 0x3D, 0x1C, 0x72, 0x3C, 0x0A, 0x41, 0x5E, 0x0E,
	0x1A, 0x55, 0x1B, 0x33, 0x24, 0x08, 0x0B, 0x16, 0x18, 0x34, 0x27, 0x0F,
	0x58, 0x5C, 0x20, 0x3E, 0x2D, 0x01, 0x5D, 0x29, 0x5D, 0x4E, 0x0A, 0x01,
	0x71, 0x09, 0x19, 0x0C, 0x52, 0x75, 0x1A, 0x4E, 0x58, 0x24, 0x24, 0x36,
	0x12, 0x20, 0x03, 0x04, 0x39, 0x57, 0x02, 0x07, 0x08, 0x43, 0x2D, 0x5A,
	0x3D, 0x2D, 0x25, 0x2F, 0x5C, 0x5E, 0x75, 0x43, 0x56, 0x28, 0x06, 0x6D,
	0x09, 0x02, 0x3E, 0x27, 0x77, 0x2E, 0x08, 0x1A, 0x39, 0x77, 0x35, 0x59,
	0x02, 0x59, 0x2F, 0x0A, 0x16, 0x1B, 0x27, 0x2B, 0x1E, 0x11, 0x08, 0x08,
	0x7B, 0x2F, 0x23, 0x41, 0x1B, 0x12, 0x0A, 0x0E, 0x09, 0x3E, 0x77, 0x5B,
	0x15, 0x34, 0x00, 0x33, 0x5A, 0x35, 0x5B, 0x5C, 0x11, 0x43, 0x33, 0x17,
	0x12, 0x34, 0x5B, 0x06, 0x04, 0x52, 0x2B, 0x23, 0x37, 0x19, 0x0A, 0x71,
	0x5B, 0x25, 0x34, 0x52, 0x34, 0x02, 0x57, 0x59, 0x08, 0x1B, 0x43, 0x28,
	0x08, 0x06, 0x26, 0x3C, 0x22, 0x18, 0x19, 0x24, 0x0A, 0x17, 0x36, 0x0C,
	0x2F, 0x5E, 0x32, 0x0A, 0x5C, 0x33, 0x3D, 0x1B, 0x19, 0x3C, 0x16, 0x5B,
	0x35, 0x0C, 0x0E, 0x20, 0x0A, 0x17, 0x03, 0x13, 0x33, 0x36, 0x14, 0x1A,
	0x1A, 0x24, 0x09, 0x57, 0x1F, 0x12, 0x1A, 0x0E, 0x10, 0x0C, 0x29, 0x69,
	0x38, 0x35, 0x34, 0x2E, 0x70, 0x0F, 0x4E, 0x05, 0x39, 0x70, 0x14, 0x30,
	0x5D, 0x40, 0x34, 0x08, 0x58, 0x14, 0x24, 0x77, 0x55, 0x14, 0x5B, 0x5D,
	0x2B, 0x5C, 0x20, 0x1C, 0x1D, 0x20, 0x5B, 0x26, 0x08, 0x08, 0x75, 0x14,
	0x2F, 0x3C, 0x1B, 0x05, 0x07, 0x3B, 0x5B, 0x1A, 0x7B, 0x15, 0x56, 0x5B,
	0x5A, 0x2E, 0x1A, 0x07, 0x20, 0x19, 0x28, 0x0A, 0x50, 0x05, 0x0D, 0x23,
	0x07, 0x59, 0x5B, 0x3A, 0x24, 0x5F, 0x34, 0x21, 0x1E, 0x33, 0x39, 0x54,
	0x34, 0x2E, 0x30, 0x25, 0x58, 0x37, 0x0A, 0x38, 0x02, 0x0C, 0x18, 0x06,
	0x74, 0x3A, 0x28, 0x0C, 0x59, 0x69, 0x1F, 0x58, 0x39, 0x2F, 0x23, 0x55,
	0x57, 0x56, 0x59, 0x05, 0x0D, 0x4A, 0x1A, 0x25, 0x74, 0x0E, 0x28, 0x5B,
	0x07, 0x26, 0x14, 0x00, 0x08, 0x44, 0x71, 0x15, 0x34, 0x19, 0x59, 0x36,
	0x59, 0x4A, 0x5A, 0x13, 0x7A, 0x02, 0x36, 0x08, 0x40, 0x27, 0x1B, 0x23,
	0x20, 0x0A, 0x36, 0x1B, 0x56, 0x58, 0x3B, 0x0E, 0x01, 0x36, 0x29, 0x31,
	0x24, 0x3C, 0x53, 0x22, 0x05, 0x24, 0x38, 0x22, 0x39, 0x07, 0x03, 0x2A,
	0x16, 0x09, 0x5E, 0x6D, 0x09, 0x23, 0x58, 0x5E, 0x26, 0x08, 0x08, 0x17,
	0x44, 0x0F, 0x0E, 0x29, 0x0C, 0x06, 0x36, 0x24, 0x51, 0x5A, 0x53, 0x33,
	0x18, 0x08, 0x34, 0x00, 0x38, 0x47, 0x56, 0x07, 0x0E, 0x72, 0x02, 0x2A,
	0x59, 0x5B, 0x7B, 0x1D, 0x2A, 0x57, 0x5A, 0x28, 0x1B, 0x12, 0x45, 0x29,
	0x0C, 0x5E, 0x2E, 0x19, 0x03, 0x10, 0x20, 0x36, 0x16, 0x26, 0x2C, 0x06,
	0x55, 0x2F, 0x08, 0x06, 0x54, 0x36, 0x21, 0x3B, 0x27, 0x28, 0x26, 0x41,
	0x40, 0x10, 0x2F, 0x53, 0x3F, 0x19, 0x25, 0x25, 0x55, 0x3D, 0x5B, 0x07,
	0x25, 0x59, 0x07, 0x2A, 0x06, 0x15, 0x26, 0x3F, 0x1A, 0x0E, 0x1D, 0x0F,
	0x24, 0x33, 0x7B, 0x3C, 0x51, 0x5A, 0x3F, 0x00, 0x2E, 0x06, 0x19, 0x1E,
	0x17, 0x55, 0x10, 0x0F, 0x20, 0x05, 0x5C, 0x37, 0x3D, 0x03, 0x36, 0x47,
	0x17, 0x27, 0x1B, 0x7B, 0x0B, 0x51, 0x17, 0x40, 0x6D, 0x06, 0x2F, 0x1F,
	0x27, 0x24, 0x3A, 0x0D, 0x5E, 0x39, 0x35, 0x08, 0x54, 0x00, 0x18, 0x27,
	0x3D, 0x30, 0x04, 0x52, 0x06, 0x29, 0x35, 0x34, 0x32, 0x76, 0x25, 0x10,
	0x39, 0x5B, 0x2E, 0x55, 0x54, 0x0B, 0x1F, 0x04, 0x15, 0x1B, 0x3F, 0x1A,
	0x71, 0x2B, 0x0F, 0x5A, 0x0F, 0x2E, 0x19, 0x26, 0x3E, 0x5A, 0x75, 0x3E,
	0x2E, 0x2C, 0x19, 0x2B, 0x01, 0x35, 0x24, 0x59, 0x7A, 0x04, 0x06, 0x5E,
	0x3D, 0x6D, 0x27, 0x07, 0x0F, 0x59, 0x35, 0x1F, 0x17, 0x3D, 0x04, 0x05,
	0x1A, 0x35, 0x16, 0x3F, 0x21, 0x1C, 0x32, 0x2B, 0x0D, 0x2E, 0x5D, 0x38,
	0x18, 0x03, 0x23, 0x36, 0x33, 0x3F, 0x32, 0x34, 0x3C, 0x08, 0x5E, 0x1A,
	0x08, 0x3F, 0x2F, 0x24, 0x27, 0x04, 0x18, 0x0F, 0x3F, 0x19, 0x18, 0x19,
	0x27, 0x18, 0x5A, 0x2D, 0x27, 0x17, 0x1A, 0x52, 0x77, 0x01, 0x22, 0x16,
	0x39, 0x07, 0x15, 0x17, 0x56, 0x53, 0x04, 0x08, 0x25, 0x2F, 0x1A, 0x34,
	0x0E, 0x59, 0x2C, 0x31, 0x6D, 0x0F, 0x0D, 0x25, 0x1F, 0x36, 0x05, 0x37,
	0x59, 0x2C, 0x71, 0x02, 0x11, 0x20, 0x02, 0x70, 0x16, 0x0B, 0x1C, 0x0A,
	0x03, 0x3A, 0x27, 0x34, 0x0E, 0x0F, 0x07, 0x22, 0x45, 0x18, 0x14, 0x00,
	0x54, 0x00, 0x5A, 0x2E, 0x1A, 0x28, 0x27, 0x29, 0x34, 0x34, 0x10, 0x22,
	0x21, 0x00, 0x39, 0x17, 0x37, 0x02, 0x14, 0x23, 0x0E, 0x5B, 0x08, 0x0F,
	0x3F, 0x55, 0x05, 0x39, 0x14, 0x54, 0x17, 0x36, 0x29, 0x3B, 0x27, 0x2A,
	0x5E, 0x52, 0x2B, 0x59, 0x18, 0x1A, 0x52, 0x27, 0x06, 0x0A, 0x5F, 0x27,
	0x32, 0x08, 0x58, 0x1F, 0x07, 0x15, 0x3B, 0x12, 0x56, 0x11, 0x7B, 0x0B,
	0x0F, 0x3A, 0x23, 0x74, 0x28, 0x36, 0x5A, 0x00, 0x25, 0x38, 0x4A, 0x24,
	0x2E, 0x01, 0x07, 0x2D, 0x1E, 0x0A, 0x10, 0x27, 0x59, 0x0F, 0x1F, 0x2B,
	0x07, 0x28, 0x5F, 0x23, 0x10, 0x1E, 0x2B, 0x2B, 0x0E, 0x1A, 0x29, 0x2E,
	0x26, 0x39, 0x11, 0x2F, 0x27, 0x5E, 0x1F, 0x0E, 0x38, 0x55, 0x3C, 0x02,
	0x76, 0x16, 0x39, 0x2F, 0x53, 0x0C, 0x1A, 0x0F, 0x14, 0x18, 0x3B, 0x3F,
	0x26, 0x2A, 0x1B, 0x0B, 0x2E, 0x18, 0x27, 0x20, 0x7A, 0x0F, 0x14, 0x57,
	0x26, 0x24, 0x38, 0x08, 0x0C, 0x53, 0x35, 0x1D, 0x25, 0x5F, 0x0C, 0x17,
	0x35, 0x05, 0x41, 0x02, 0x00, 0x35, 0x24, 0x09, 0x29, 0x18, 0x58, 0x37,
	0x36, 0x02, 0x29, 0x1E, 0x2F, 0x3D, 0x5B, 0x33, 0x20, 0x00, 0x1D, 0x1F,
	0x7A, 0x1D, 0x2D, 0x36, 0x3A, 0x77, 0x25, 0x15, 0x3A, 0x02, 0x14, 0x04,
	0x2D, 0x3D, 0x1D, 0x00, 0x05, 0x30, 0x04, 0x31, 0x3A, 0x27, 0x32, 0x03,
	0x1B, 0x1B, 0x29, 0x05, 0x34, 0x06, 0x1B, 0x54, 0x38, 0x3B, 0x21, 0x33,
	0x2E, 0x08, 0x58, 0x28, 0x20, 0x21, 0x24, 0x08, 0x3C, 0x23, 0x35, 0x4A,
	0x0C, 0x28, 0x7B, 0x2E, 0x13, 0x07, 0x2C, 0x32, 0x39, 0x17, 0x37, 0x19,
	0x7A, 0x3F, 0x19, 0x20, 0x19, 0x38, 0x3D, 0x19, 0x3B, 0x40, 0x36, 0x35,
	0x25, 0x14, 0x31, 0x2F, 0x5D, 0x30, 0x07, 0x53, 0x3A, 0x29, 0x34, 0x0D,
	0x59, 0x3A, 0x36, 0x0E, 0x37, 0x44, 0x13, 0x1D, 0x30, 0x0F, 0x13, 0x14,
	0x16, 0x26, 0x06, 0x52, 0x0D, 0x0B, 0x26, 0x56, 0x01, 0x3A, 0x19, 0x09,
	0x02, 0x31, 0x16, 0x23, 0x08, 0x29, 0x00, 0x76, 0x2B, 0x05, 0x2C, 0x1C,
	0x29, 0x20, 0x00, 0x28, 0x39, 0x0E, 0x2B, 0x31, 0x36, 0x5E, 0x70, 0x1A,
	0x04, 0x1F, 0x53, 0x24, 0x26, 0x16, 0x2D, 0x07, 0x2D, 0x04, 0x14, 0x0B,
	0x28, 0x0E, 0x47, 0x0E, 0x22, 0x20, 0x09, 0x1E, 0x06, 0x3A, 0x2C, 0x37,
	0x04, 0x08, 0x23, 0x53, 0x71, 0x5C, 0x25, 0x5D, 0x04, 0x07, 0x2F, 0x09,
	0x1C, 0x11, 0x06, 0x29, 0x2C, 0x14, 0x28, 0x29, 0x00, 0x11, 0x25, 0x5C,
	0x72, 0x39, 0x39, 0x2C, 0x19, 0x75, 0x08, 0x0F, 0x1E, 0x22, 0x36, 0x14,
	0x08, 0x3F, 0x32, 0x2C, 0x1C, 0x12, 0x3C, 0x0A, 0x7A, 0x0E, 0x15, 0x22,
	0x1B, 0x05, 0x07, 0x55, 0x27, 0x0E, 0x31, 0x23, 0x52, 0x38, 0x25, 0x35,
	0x27, 0x51, 0x5C, 0x12, 0x36, 0x19, 0x4A, 0x0B, 0x00, 0x10, 0x26, 0x0B,
	0x5C, 0x52, 0x1B, 0x0D, 0x53, 0x17, 0x31, 0x09, 0x38, 0x2B, 0x26, 0x07,
	0x1B, 0x22, 0x53, 0x25, 0x33, 0x2C, 0x0F, 0x10, 0x36, 0x31, 0x13, 0x19,
	0x0D, 0x02, 0x1A, 0x71, 0x3F, 0x0E, 0x5E, 0x0E, 0x00, 0x2E, 0x34, 0x09,
	0x08, 0x35, 0x59, 0x05, 0x38, 0x52, 0x23, 0x15, 0x09, 0x1D, 0x27, 0x17,
	0x5E, 0x58, 0x2F, 0x5F, 0x34, 0x2F, 0x10, 0x09, 0x0D, 0x01, 0x29, 0x04,
	0x0B, 0x04, 0x29, 0x03, 0x02, 0x5D, 0x25, 0x17, 0x18, 0x33, 0x2F, 0x0C,
	0x24, 0x36, 0x33, 0x45, 0x05, 0x26, 0x35, 0x02, 0x0B, 0x19, 0x0D, 0x27,
	0x58, 0x59, 0x27, 0x75, 0x09, 0x32, 0x39, 0x07, 0x72, 0x1F, 0x17, 0x1A,
	0x1B, 0x17, 0x2E, 0x17, 0x1E, 0x25, 0x69, 0x5C, 0x0E, 0x57, 0x44, 0x31,
	0x22, 0x35, 0x23, 0x09, 0x0B, 0x24, 0x14, 0x1A, 0x18, 0x26, 0x03, 0x03,
	0x04, 0x0D, 0x10, 0x1E, 0x0B, 0x59, 0x3D, 0x04, 0x3D, 0x0C, 0x2B, 0x53,
	0x11, 0x3A, 0x33, 0x25, 0x32, 0x2D, 0x1B, 0x1B, 0x2A, 0x1C, 0x71, 0x2A,
	0x00, 0x5E, 0x53, 0x29, 0x0B, 0x22, 0x2C, 0x59, 0x74, 0x18, 0x18, 0x16,
	0x3A, 0x77, 0x0F, 0x2E, 0x56, 0x1D, 0x20, 0x5C, 0x29, 0x59, 0x5E, 0x24,
	0x02, 0x11, 0x5A, 0x39, 0x06, 0x39, 0x36, 0x19, 0x3A, 0x36, 0x35, 0x59,
	0x5F, 0x2D, 0x20, 0x47, 0x58, 0x03, 0x2A, 0x72, 0x34, 0x15, 0x23, 0x2E,
	0x00, 0x1C, 0x55, 0x05, 0x08, 0x17, 0x1C, 0x52, 0x5F, 0x2D, 0x20, 0x2A,
	0x2E, 0x05, 0x06, 0x33, 0x5D, 0x0C, 0x5D, 0x5D, 0x32, 0x47, 0x14, 0x00,
	0x12, 0x16, 0x08, 0x22, 0x58, 0x31, 0x7B, 0x05, 0x11, 0x38, 0x31, 0x2F,
	0x21, 0x50, 0x3C, 0x28, 0x0E, 0x3F, 0x36, 0x3B, 0x19, 0x3B, 0x21, 0x06,
	0x2A, 0x53, 0x30, 0x06, 0x14, 0x19, 0x06, 0x1A, 0x43, 0x59, 0x08, 0x05,
	0x07, 0x43, 0x0D, 0x59, 0x26, 0x12, 0x20, 0x52, 0x0A, 0x1E, 0x16, 0x02,
	0x35, 0x0D, 0x3D, 0x75, 0x21, 0x22, 0x58, 0x12, 0x26, 0x39, 0x36, 0x5F,
	0x2C, 0x01, 0x16, 0x37, 0x05, 0x1A, 0x07, 0x38, 0x39, 0x5A, 0x3B, 0x38,
	0x54, 0x29, 0x0B, 0x24, 0x18, 0x0F, 0x52, 0x1C, 0x0D, 0x30, 0x1D, 0x0C,
	0x16, 0x3C, 0x24, 0x3D, 0x00, 0x5A, 0x5C, 0x07, 0x1C, 0x08, 0x34, 0x23,
	0x08, 0x38, 0x28, 0x1A, 0x0C, 0x15, 0x0A, 0x0D, 0x2B, 0x39, 0x16, 0x0B,
	0x57, 0x06, 0x1D, 0x1B, 0x18, 0x14, 0x01, 0x1C, 0x1A, 0x1E, 0x12, 0x04,
	0x2A, 0x71, 0x1C, 0x36, 0x01, 0x01, 0x11, 0x20, 0x3B, 0x17, 0x33, 0x72,
	0x55, 0x30, 0x58, 0x3E, 0x0E, 0x3E, 0x04, 0x28, 0x0C, 0x2A, 0x04, 0x0F,
	0x23, 0x12, 0x6D, 0x15, 0x2C, 0x1A, 0x2C, 0x06, 0x1B, 0x0B, 0x17, 0x2F,
	0x34, 0x0A, 0x18, 0x2A, 0x1C, 0x36, 0x1F, 0x08, 0x09, 0x3C, 0x3A, 0x29,
	0x54, 0x2D, 0x3C, 0x2E, 0x1C, 0x10, 0x08, 0x01, 0x11, 0x1F, 0x04, 0x22,
	0x29, 0x11, 0x38, 0x26, 0x24, 0x08, 0x20, 0x0B, 0x20, 0x34, 0x52, 0x2C,
	0x26, 0x07, 0x2F, 0x3B, 0x07, 0x0B, 0x13, 0x1E, 0x07, 0x05, 0x3E, 0x25,
	0x3A, 0x08, 0x73, 0x0D, 0x28, 0x3F, 0x04, 0x36, 0x5C, 0x24, 0x1D, 0x3A,
	0x0F, 0x54, 0x50, 0x2D, 0x44, 0x37, 0x26, 0x0E, 0x21, 0x05, 0x76, 0x55,
	0x29, 0x00, 0x0E, 0x21, 0x0D, 0x29, 0x19, 0x2E, 0x34, 0x5D, 0x11, 0x25,
	0x25, 0x38, 0x01, 0x04, 0x38, 0x3C, 0x2B, 0x0B, 0x09, 0x57, 0x12, 0x09,
	0x39, 0x26, 0x37, 0x5A, 0x0A, 0x08, 0x0D, 0x1C, 0x5C, 0x71, 0x05, 0x25,
	0x2A, 0x04, 0x31, 0x34, 0x26, 0x05, 0x05, 0x06, 0x20, 0x16, 0x1A, 0x09,
	0x72, 0x2E, 0x52, 0x08, 0x22, 0x36, 0x5F, 0x2A, 0x27, 0x1F, 0x74, 0x0D,
	0x3B, 0x16, 0x23, 0x24, 0x00, 0x12, 0x0B, 0x11, 0x11, 0x04, 0x2F, 0x22,
	0x03, 0x72, 0x35, 0x0D, 0x0A, 0x32, 0x21, 0x08, 0x00, 0x2D, 0x1A, 0x0C,
	0x35, 0x0F, 0x41, 0x40, 0x12, 0x2E, 0x03, 0x14, 0x53, 0x69, 0x0F, 0x0D,
	0x2D, 0x23, 0x21, 0x04, 0x00, 0x23, 0x3B, 0x69, 0x22, 0x59, 0x2C, 0x33,
	0x07, 0x2D, 0x2D, 0x2F, 0x27, 0x77, 0x07, 0x53, 0x03, 0x31, 0x72, 0x08,
	0x04, 0x29, 0x07, 0x35, 0x3B, 0x10, 0x2C, 0x33, 0x35, 0x25, 0x32, 0x0B,
	0x05, 0x08, 0x29, 0x0C, 0x02, 0x0C, 0x70, 0x20, 0x4A, 0x3E, 0x12, 0x0E,
	0x34, 0x52, 0x0C, 0x2D, 0x0B, 0x15, 0x27, 0x0B, 0x11, 0x01, 0x39, 0x0D,
	0x28, 0x09, 0x32, 0x2A, 0x37, 0x22, 0x11, 0x1B, 0x04, 0x09, 0x02, 0x07,
	0x07, 0x35, 0x4E, 0x0C, 0x5F, 0x32, 0x00, 0x09, 0x2F, 0x21, 0x69, 0x07,
	0x2D, 0x38, 0x03, 0x0E, 0x47, 0x24, 0x3B, 0x1B, 0x17, 0x1C, 0x29, 0x36,
	0x06, 0x3B, 0x25, 0x04, 0x0A, 0x1C, 0x72, 0x18, 0x53, 0x36, 0x02, 0x01,
	0x3A, 0x4E, 0x0C, 0x2A, 0x01, 0x5F, 0x12, 0x23, 0x1C, 0x71, 0x1E, 0x18,
	0x1D, 0x00, 0x34, 0x3F, 0x19, 0x3C, 0x06, 0x3A, 0x1D, 0x04, 0x2F, 0x02,
	0x3A, 0x08, 0x0A, 0x3B, 0x19, 0x69, 0x5A, 0x32, 0x2D, 0x06, 0x21, 0x01,
	0x0F, 0x00, 0x1C, 0x1B, 0x1F, 0x28, 0x07, 0x3D, 0x0E, 0x5F, 0x15, 0x3B,
	0x31, 0x38, 0x15, 0x59, 0x59, 0x22, 0x0C, 0x1F, 0x03, 0x25, 0x5C, 0x11,
	0x14, 0x58, 0x37, 0x28, 0x1A, 0x3A, 0x53, 0x34, 0x3C, 0x13, 0x01, 0x35,
	0x1D, 0x5B, 0x11, 0x3F, 0x27, 0x27, 0x44, 0x13, 0x39, 0x15, 0x03, 0x1A,
	0x27, 0x18, 0x00, 0x56, 0x19, 0x07, 0x3E, 0x19, 0x2B, 0x01, 0x73, 0x26,
	0x16, 0x3B, 0x18, 0x09, 0x5C, 0x22, 0x18, 0x0F, 0x03, 0x2F, 0x50, 0x3E,
	0x24, 0x06, 0x1E, 0x0D, 0x5B, 0x5B, 0x69, 0x1D, 0x09, 0x07, 0x2F, 0x2C,
	0x08, 0x33, 0x06, 0x5E, 0x13, 0x5B, 0x2B, 0x1D, 0x33, 0x14, 0x59, 0x54,
	0x22, 0x08, 0x25, 0x0D, 0x0E, 0x05, 0x33, 0x14, 0x1B, 0x0F, 0x00, 0x26,
	0x36, 0x1D, 0x20, 0x28, 0x52, 0x71, 0x18, 0x56, 0x1E, 0x3E, 0x30, 0x5B,
	0x22, 0x0D, 0x23, 0x21, 0x0A, 0x11, 0x22, 0x3A, 0x2E, 0x24, 0x15, 0x0D,
	0x1A, 0x30, 0x38, 0x17, 0x3B, 0x1B, 0x69, 0x5B, 0x2D, 0x5F, 0x2E, 0x74,
	0x02, 0x10, 0x0B, 0x5B, 0x12, 0x5C, 0x0D, 0x1E, 0x58, 0x72, 0x07, 0x11,
	0x18, 0x1B, 0x1A, 0x3F, 0x07, 0x02, 0x5F, 0x38, 0x5B, 0x0F, 0x58, 0x03,
	0x29, 0x1E, 0x50, 0x5B, 0x38, 0x34, 0x1A, 0x25, 0x02, 0x3B, 0x0F, 0x5F,
	0x55, 0x1B, 0x5E, 0x6D, 0x39, 0x15, 0x1C, 0x05, 0x01, 0x0E, 0x0B, 0x02,
	0x1F, 0x14, 0x20, 0x00, 0x57, 0x5A, 0x05, 0x15, 0x2B, 0x5F, 0x20, 0x77,
	0x43, 0x24, 0x1C, 0x40, 0x76, 0x05, 0x17, 0x1E, 0x1E, 0x3B, 0x05, 0x0D,
	0x1A, 0x5B, 0x12, 0x26, 0x52, 0x06, 0x20, 0x2E, 0x43, 0x37, 0x07, 0x07,
	0x7B, 0x24, 0x2A, 0x38, 0x01, 0x2F, 0x0F, 0x13, 0x5B, 0x3D, 0x69, 0x1D,
	0x37, 0x24, 0x5E, 0x0B, 0x1C, 0x07, 0x16, 0x33, 0x09, 0x3E, 0x52, 0x3E,
	0x3E, 0x17, 0x1C, 0x17, 0x05, 0x1F, 0x0B, 0x47, 0x2D, 0x5E, 0x2C, 0x32,
	0x3C, 0x24, 0x1C, 0x5C, 0x32, 0x39, 0x13, 0x1C, 0x38, 0x17, 0x08, 0x04,
	0x1F, 0x05, 0x34, 0x43, 0x59, 0x3F, 0x23, 0x37, 0x1A, 0x0C, 0x28, 0x28,
	0x36, 0x34, 0x26, 0x37, 0x59, 0x7B, 0x5A, 0x34, 0x04, 0x00, 0x37, 0x0E,
	0x02, 0x1D, 0x0D, 0x3A, 0x2F, 0x08, 0x5D, 0x1E, 0x6D, 0x05, 0x26, 0x02,
	0x44, 0x15, 0x22, 0x2A, 0x45, 0x5D, 0x27, 0x39, 0x58, 0x1E, 0x2C, 0x2A,
	0x39, 0x0F, 0x03, 0x5A, 0x37, 0x0F, 0x07, 0x22, 0x07, 0x24, 0x0E, 0x2D,
	0x02, 0x3B, 0x23, 0x3E, 0x51, 0x00, 0x05, 0x04, 0x39, 0x26, 0x00, 0x0D,
	0x10, 0x2B, 0x0F, 0x08, 0x38, 0x2F, 0x01, 0x4E, 0x3A, 0x26, 0x2F, 0x09,
	0x32, 0x25, 0x33, 0x74, 0x27, 0x37, 0x39, 0x12, 0x30, 0x5D, 0x32, 0x2A,
	0x1A, 0x77, 0x47, 0x0F, 0x0A, 0x2F, 0x3A, 0x3F, 0x4A, 0x0C, 0x01, 0x11,
	0x3C, 0x0A, 0x56, 0x1B, 0x24, 0x0D, 0x32, 0x5E, 0x5C, 0x74, 0x27, 0x51,
	0x36, 0x5D, 0x05, 0x39, 0x07, 0x1C, 0x09, 0x11, 0x54, 0x36, 0x17, 0x07,
	0x7B, 0x26, 0x27, 0x3D, 0x0D, 0x10, 0x07, 0x10, 0x45, 0x32, 0x36, 0x02,
	0x1B, 0x14, 0x59, 0x27, 0x5D, 0x51, 0x34, 0x1B, 0x24, 0x34, 0x20, 0x02,
	0x0D, 0x73, 0x3F, 0x38, 0x0D, 0x25, 0x36, 0x28, 0x11, 0x38, 0x27, 0x69,
	0x5B, 0x54, 0x3A, 0x59, 0x34, 0x08, 0x52, 0x0A, 0x05, 0x1A, 0x00, 0x36,
	0x0D, 0x29, 0x20, 0x15, 0x25, 0x1C, 0x08, 0x08, 0x04, 0x56, 0x3E, 0x3A,
	0x0F, 0x27, 0x07, 0x21, 0x04, 0x31, 0x58, 0x2E, 0x20, 0x03, 0x29, 0x14,
	0x00, 0x38, 0x22, 0x20, 0x1A, 0x20, 0x2A, 0x1F, 0x0F, 0x28, 0x0B, 0x3A,
	0x21, 0x0F, 0x2D, 0x24, 0x20, 0x28, 0x0F, 0x3E, 0x1B, 0x1E, 0x01, 0x10,
	0x3B, 0x35, 0x19, 0x58, 0x2F, 0x3C, 0x55, 0x00, 0x38, 0x0A, 0x00, 0x22,
	0x1B, 0x2A, 0x01, 0x28, 0x30, 0x0C, 0x53, 0x36, 0x1E, 0x55, 0x21, 0x52,
	0x30, 0x0E, 0x51, 0x1A, 0x44, 0x71, 0x08, 0x57, 0x18, 0x52, 0x12, 0x5B,
	0x0F, 0x0A, 0x5C, 0x34, 0x55, 0x29, 0x58, 0x05, 0x7B, 0x16, 0x14, 0x57,
	0x58, 0x69, 0x02, 0x58, 0x3A, 0x1E, 0x7B, 0x5F, 0x04, 0x1C, 0x44, 0x16,
	0x47, 0x52, 0x08, 0x38, 0x69, 0x5B, 0x52, 0x57, 0x58, 0x34, 0x59, 0x29,
	0x0C, 0x5F, 0x1B, 0x25, 0x2F, 0x0F, 0x31, 0x34, 0x5B, 0x0D, 0x27, 0x5B,
	0x0E, 0x06, 0x2D, 0x2B, 0x52, 0x71, 0x35, 0x11, 0x29, 0x01, 0x7A, 0x35,
	0x55, 0x1A, 0x53, 0x00, 0x27, 0x33, 0x01, 0x1F, 0x28, 0x3C, 0x23, 0x18,
	0x09, 0x00, 0x3F, 0x2F, 0x27, 0x39, 0x03, 0x54, 0x30, 0x23, 0x09, 0x76,
	0x36, 0x16, 0x21, 0x5F, 0x00, 0x2D, 0x30, 0x34, 0x5F, 0x7B, 0x3F, 0x26,
	0x0D, 0x27, 0x72, 0x23, 0x2C, 0x1D, 0x31, 0x06, 0x28, 0x07, 0x28, 0x25,
	0x1B, 0x25, 0x13, 0x29, 0x04, 0x76, 0x5C, 0x30, 0x03, 0x0C, 0x1B, 0x15,
	0x19, 0x09, 0x53, 0x13, 0x2A, 0x14, 0x2C, 0x0D, 0x12, 0x3E, 0x12, 0x04,
	0x39, 0x07, 0x2E, 0x38, 0x2C, 0x09, 0x0B, 0x04, 0x0E, 0x2A, 0x2C, 0x07,
	0x3D, 0x11, 0x2C, 0x5E, 0x25, 0x29, 0x02, 0x06, 0x19, 0x03, 0x23, 0x54,
	0x2A, 0x2D, 0x06, 0x0A, 0x23, 0x25, 0x2E, 0x7B, 0x3B, 0x20, 0x08, 0x3A,
	0x70, 0x2D, 0x32, 0x18, 0x38, 0x35, 0x21, 0x57, 0x09, 0x2C, 0x1B, 0x3D,
	0x35, 0x01, 0x23, 0x0F, 0x2E, 0x1B, 0x19, 0x2F, 0x2D, 0x3D, 0x1B, 0x1C,
	0x2A, 0x73, 0x58, 0x16, 0x19, 0x09, 0x7B, 0x16, 0x34, 0x18, 0x0C, 0x74,
	0x29, 0x13, 0x5C, 0x28, 0x17, 0x2D, 0x54, 0x17, 0x21, 0x23, 0x2E, 0x53,
	0x2B, 0x5F, 0x10, 0x19, 0x55, 0x26, 0x3A, 0x03, 0x06, 0x32, 0x28, 0x3E,
	0x76, 0x24, 0x30, 0x2F, 0x1E, 0x72, 0x2F, 0x55, 0x2A, 0x5C, 0x0B, 0x20,
	0x0E, 0x2A, 0x1E, 0x07, 0x14, 0x18, 0x2F, 0x27, 0x03, 0x29, 0x2C, 0x09,
	0x3B, 0x03, 0x0F, 0x54, 0x2B, 0x01, 0x03, 0x2B, 0x30, 0x07, 0x33, 0x0B,
	0x29, 0x12, 0x2A, 0x21, 0x07, 0x22, 0x57, 0x2C, 0x05, 0x03, 0x21, 0x55,
	0x2C, 0x53, 0x0B, 0x02, 0x0A, 0x3E, 0x26, 0x03, 0x22, 0x51, 0x26, 0x5F,
	0x00, 0x02, 0x28, 0x1E, 0x5F, 0x01, 0x2B, 0x59, 0x5C, 0x29, 0x26, 0x2E,
	0x55, 0x0C, 0x3C, 0x34, 0x5C, 0x23, 0x23, 0x22, 0x23, 0x05, 0x23, 0x36,
	0x2A, 0x30, 0x5A, 0x27, 0x01, 0x22, 0x17, 0x34, 0x53, 0x39, 0x1E, 0x09,
	0x39, 0x23, 0x23, 0x22, 0x27, 0x05, 0x25, 0x14, 0x2A, 0x04, 0x18, 0x23,
	0x23, 0x2A, 0x11, 0x36, 0x25, 0x45, 0x0C, 0x0E, 0x03, 0x30, 0x26, 0x22,
	0x03, 0x07, 0x20, 0x06, 0x29, 0x00, 0x23, 0x30, 0x27, 0x1C, 0x0A, 0x1E,
	0x0C, 0x3D, 0x27, 0x17, 0x28, 0x26, 0x3C, 0x2F, 0x35, 0x21, 0x56, 0x20,
	0x2E, 0x20, 0x25, 0x22, 0x5C, 0x0A, 0x17, 0x59, 0x17, 0x04, 0x40, 0x07,
	0x07, 0x23, 0x3E, 0x22, 0x27, 0x35, 0x23, 0x24, 0x27, 0x10, 0x24, 0x18,
	0x2C, 0x5A, 0x29, 0x2F, 0x14, 0x24, 0x06, 0x0A, 0x07, 0x20, 0x2A, 0x00,
	0x17, 0x1F, 0x20, 0x36, 0x31, 0x25, 0x06, 0x50, 0x16, 0x11, 0x1B, 0x2D,
	0x08, 0x1D, 0x12, 0x2A, 0x1A, 0x0F, 0x2D, 0x0A, 0x25, 0x26, 0x02, 0x06,
	0x38, 0x07, 0x2B, 0x14, 0x23, 0x20, 0x24, 0x34, 0x58, 0x3B, 0x22, 0x28,
	0x3D, 0x02, 0x0F, 0x04, 0x73, 0x14, 0x10, 0x06, 0x38, 0x16, 0x0B, 0x17,
	0x19, 0x28, 0x70, 0x18, 0x59, 0x0F, 0x04, 0x32, 0x07, 0x20, 0x59, 0x0C,
	0x1B, 0x3D, 0x17, 0x27, 0x2F, 0x77, 0x0F, 0x2D, 0x0D, 0x20, 0x7A, 0x00,
	0x30, 0x05, 0x18, 0x35, 0x28, 0x4A, 0x06, 0x03, 0x00, 0x34, 0x36, 0x26,
	0x09, 0x13, 0x0D, 0x2C, 0x0C, 0x0C, 0x36, 0x14, 0x12, 0x2F, 0x59, 0x03,
	0x5A, 0x04, 0x5D, 0x2A, 0x04, 0x15, 0x23, 0x00, 0x2A, 0x35, 0x0D, 0x50,
	0x06, 0x5C, 0x30, 0x28, 0x2E, 0x01, 0x2F, 0x7B, 0x1E, 0x00, 0x26, 0x1E,
	0x31, 0x2D, 0x53, 0x2F, 0x3C, 0x16, 0x36, 0x30, 0x3C, 0x5A, 0x25, 0x24,
	0x12, 0x25, 0x00, 0x36, 0x47, 0x23, 0x41, 0x5C, 0x00, 0x24, 0x22, 0x1A,
	0x23, 0x24, 0x0B, 0x07, 0x5B, 0x29, 0x0E, 0x2D, 0x2F, 0x2C, 0x03, 0x12,
	0x1A, 0x53, 0x2B, 0x0F, 0x35, 0x2E, 0x2C, 0x0A, 0x1C, 0x04, 0x0F, 0x0A,
	0x5C, 0x2A, 0x03, 0x03, 0x15, 0x3F, 0x0D, 0x6D, 0x0B, 0x2B, 0x19, 0x25,
	0x27, 0x27, 0x16, 0x04, 0x3A, 0x33, 0x5C, 0x19, 0x2A, 0x12, 0x2A, 0x5C,
	0x30, 0x27, 0x0C, 0x12, 0x0F, 0x08, 0x3A, 0x0C, 0x2E, 0x29, 0x55, 0x27,
	0x0F, 0x13, 0x21, 0x54, 0x2C, 0x58, 0x03, 0x19, 0x23, 0x2F, 0x40, 0x13,
	0x54, 0x16, 0x2A, 0x52, 0x0D, 0x15, 0x31, 0x05, 0x2A, 0x75, 0x25, 0x20,
	0x56, 0x20, 0x29, 0x06, 0x50, 0x2A, 0x0D, 0x0B, 0x00, 0x38, 0x2D, 0x1D,
	0x27, 0x05, 0x20, 0x3B, 0x02, 0x15, 0x34, 0x20, 0x5F, 0x5D, 0x76, 0x25,
	0x25, 0x3F, 0x26, 0x18, 0x19, 0x32, 0x2B, 0x5B, 0x00, 0x21, 0x28, 0x5E,
	0x05, 0x00, 0x08, 0x06, 0x34, 0x5B, 0x6D, 0x1B, 0x20, 0x56, 0x0C, 0x37,
	0x0B, 0x2C, 0x0C, 0x0E, 0x17, 0x24, 0x00, 0x3F, 0x0E, 0x1B, 0x2F, 0x1B,
	0x08, 0x29, 0x06, 0x0D, 0x06, 0x0A, 0x26, 0x0A, 0x0A, 0x2E, 0x3B, 0x3B,
	0x20, 0x3E, 0x2A, 0x00, 0x2A, 0x6D, 0x0B, 0x0E, 0x2F, 0x26, 0x33, 0x2A,
	0x3B, 0x0D, 0x2F, 0x71, 0x29, 0x2F, 0x59, 0x03, 0x0C, 0x2D, 0x31, 0x2C,
	0x25, 0x72, 0x24, 0x30, 0x08, 0x19, 0x06, 0x22, 0x06, 0x24, 0x5D, 0x7B,
	0x1B, 0x04, 0x56, 0x3E, 0x70, 0x2D, 0x31, 0x5A, 0x2F, 0x2D, 0x25, 0x2B,
	0x17, 0x28, 0x25, 0x35, 0x18, 0x07, 0x5D, 0x07, 0x09, 0x06, 0x0D, 0x5E,
	0x05, 0x5F, 0x23, 0x28, 0x0D, 0x3B, 0x0B, 0x0B, 0x17, 0x28, 0x15, 0x2D,
	0x02, 0x5C, 0x24, 0x2A, 0x34, 0x22, 0x2A, 0x05, 0x03, 0x36, 0x0E, 0x3E,
	0x03, 0x6D, 0x27, 0x20, 0x14, 0x2A, 0x24, 0x21, 0x29, 0x5A, 0x07, 0x13,
	0x20, 0x2F, 0x37, 0x29, 0x0E, 0x2E, 0x0E, 0x28, 0x3B, 0x31, 0x25, 0x18,
	0x37, 0x20, 0x12, 0x3E, 0x22, 0x2B, 0x5B, 0x03, 0x01, 0x30, 0x0D, 0x5F,
	0x18, 0x2D, 0x1B, 0x5E, 0x3A, 0x18, 0x1B, 0x0C, 0x01, 0x24, 0x17, 0x58,
	0x12, 0x2C, 0x44, 0x0A, 0x2E, 0x05, 0x3F, 0x0F, 0x28, 0x5D, 0x20, 0x1E,
	0x12, 0x0B, 0x0D, 0x20, 0x14, 0x3C, 0x18, 0x2D, 0x31, 0x56, 0x27, 0x74,
	0x0B, 0x2E, 0x0A, 0x11, 0x2D, 0x3C, 0x53, 0x2A, 0x33, 0x03, 0x24, 0x0E,
	0x23, 0x2A, 0x24, 0x1D, 0x20, 0x03, 0x3A, 0x1A, 0x3D, 0x2D, 0x3F, 0x32,
	0x20, 0x2A, 0x00, 0x04, 0x0A, 0x08, 0x15, 0x18, 0x2B, 0x06, 0x35, 0x28,
	0x2E, 0x3F, 0x08, 0x35, 0x08, 0x23, 0x38, 0x28, 0x0E, 0x05, 0x23, 0x26,
	0x2A, 0x25, 0x35, 0x37, 0x27, 0x29, 0x13, 0x2E, 0x12, 0x09, 0x2F, 0x35,
	0x47, 0x09, 0x1F, 0x2E, 0x08, 0x2F, 0x23, 0x36, 0x2A, 0x0C, 0x5B, 0x00,
	0x2A, 0x06, 0x72, 0x21, 0x18, 0x5A, 0x29, 0x6D, 0x00, 0x02, 0x27, 0x5F,
	0x03, 0x24, 0x28, 0x0B, 0x5F, 0x0D, 0x03, 0x25, 0x5A, 0x29, 0x27, 0x3D,
	0x32, 0x19, 0x28, 0x7B, 0x28, 0x51, 0x22, 0x09, 0x35, 0x24, 0x24, 0x2C,
	0x1B, 0x1B, 0x09, 0x06, 0x14, 0x5F, 0x09, 0x0F, 0x25, 0x39, 0x03, 0x77,
	0x2B, 0x04, 0x19, 0x29, 0x2F, 0x3D, 0x4E, 0x37, 0x40, 0x16, 0x0E, 0x51,
	0x25, 0x33, 0x15, 0x1B, 0x23, 0x57, 0x2F, 0x29, 0x28, 0x0E, 0x16, 0x39,
	0x0B, 0x3C, 0x2C, 0x2F, 0x58, 0x27, 0x58, 0x0B, 0x34, 0x2A, 0x70, 0x15,
	0x20, 0x22, 0x2F, 0x04, 0x25, 0x57, 0x06, 0x58, 0x38, 0x2D, 0x2F, 0x21,
	0x0C, 0x32, 0x2D, 0x29, 0x0D, 0x0C, 0x74, 0x0B, 0x51, 0x5C, 0x3B, 0x0B,
	0x2A, 0x59, 0x0D, 0x2D, 0x24, 0x2D, 0x23, 0x06, 0x23, 0x21, 0x05, 0x37,
	0x09, 0x23, 0x0D, 0x0A, 0x30, 0x2C, 0x18, 0x05, 0x23, 0x30, 0x56, 0x1C,
	0x0A, 0x54, 0x28, 0x0B, 0x00, 0x07, 0x1F, 0x20, 0x20, 0x5B, 0x0B, 0x03,
	0x23, 0x0C, 0x00, 0x17, 0x0F, 0x25, 0x45, 0x2E, 0x13, 0x15, 0x22, 0x36,
	0x2A, 0x16, 0x5A, 0x24, 0x0D, 0x2A, 0x38, 0x24, 0x23, 0x3C, 0x11, 0x3B,
	0x2A, 0x2E, 0x01, 0x0F, 0x77, 0x2B, 0x1B, 0x2F, 0x01, 0x10, 0x28, 0x2A,
	0x1D, 0x3F, 0x75, 0x0B, 0x00, 0x3F, 0x0C, 0x14, 0x3B, 0x23, 0x45, 0x1C,
	0x3A, 0x38, 0x2C, 0x37, 0x08, 0x75, 0x2D, 0x58, 0x09, 0x24, 0x29, 0x3D,
	0x2A, 0x1C, 0x2E, 0x69, 0x35, 0x2F, 0x20, 0x20, 0x23, 0x2D, 0x4A, 0x37,
	0x29, 0x75, 0x14, 0x0D, 0x3C, 0x28, 0x00, 0x28, 0x25, 0x08, 0x2A, 0x12,
	0x03, 0x28, 0x1D, 0x13, 0x25, 0x0E, 0x10, 0x2C, 0x01, 0x0E, 0x2A, 0x23,
	0x27, 0x52, 0x25, 0x24, 0x0C, 0x3F, 0x0E, 0x1B, 0x5C, 0x54, 0x06, 0x2A,
	0x0B, 0x3F, 0x23, 0x04, 0x52, 0x05, 0x04, 0x2A, 0x01, 0x2D, 0x25, 0x22,
	0x31, 0x29, 0x5F, 0x13, 0x5A, 0x27, 0x19, 0x11, 0x03, 0x0B, 0x52, 0x2A,
	0x08, 0x13, 0x2A, 0x15, 0x39, 0x03, 0x08, 0x03, 0x26, 0x1D, 0x03, 0x7A,
	0x1B, 0x27, 0x1D, 0x3A, 0x7A, 0x06, 0x20, 0x3E, 0x24, 0x0B, 0x3A, 0x29,
	0x01, 0x23, 0x17, 0x58, 0x2D, 0x07, 0x29, 0x2E, 0x38, 0x10, 0x2F, 0x0F,
	0x0B, 0x2E, 0x12, 0x2D, 0x01, 0x2F, 0x14, 0x29, 0x01, 0x2C, 0x0F, 0x0D,
	0x14, 0x23, 0x53, 0x11, 0x15, 0x2A, 0x56, 0x52, 0x25, 0x3F, 0x11, 0x19,
	0x06, 0x2D, 0x2D, 0x29, 0x0C, 0x3A, 0x28, 0x5C, 0x25, 0x1B, 0x3A, 0x3B,
	0x1B, 0x20, 0x03, 0x1B, 0x1B, 0x26, 0x12, 0x03, 0x13, 0x03, 0x34, 0x2C,
	0x06, 0x12, 0x03, 0x2D, 0x14, 0x3F, 0x3A, 0x35, 0x09, 0x09, 0x5C, 0x29,
	0x0B, 0x07, 0x22, 0x39, 0x2A, 0x07, 0x58, 0x56, 0x3A, 0x28, 0x03, 0x1C,
	0x50, 0x09, 0x2E, 0x7A, 0x2E, 0x53, 0x2B, 0x0A, 0x3B, 0x2E, 0x36, 0x2F,
	0x0D, 0x3A, 0x5C, 0x09, 0x3B, 0x28, 0x75, 0x25, 0x04, 0x37, 0x28, 0x0E,
	0x06, 0x09, 0x28, 0x04, 0x03, 0x36, 0x38, 0x2C, 0x13, 0x77, 0x1B, 0x29,
	0x0B, 0x5B, 0x06, 0x23, 0x23, 0x1B, 0x13, 0x73, 0x0B, 0x34, 0x2D, 0x23,
	0x13, 0x2E, 0x38, 0x2F, 0x39, 0x2E, 0x5C, 0x08, 0x3B, 0x2F, 0x2E, 0x23,
	0x24, 0x41, 0x2F, 0x03, 0x36, 0x30, 0x27, 0x52, 0x00, 0x5B, 0x0A, 0x23,
	0x18, 0x07, 0x21, 0x54, 0x09, 0x3F, 0x74, 0x2E, 0x56, 0x2F, 0x21, 0x76,
	0x43, 0x08, 0x1F, 0x29, 0x36, 0x20, 0x30, 0x09, 0x0D, 0x21, 0x2E, 0x53,
	0x5F, 0x53, 0x04, 0x24, 0x28, 0x3E, 0x26, 0x00, 0x20, 0x58, 0x5E, 0x00,
	0x17, 0x2B, 0x17, 0x23, 0x2A, 0x71, 0x0D, 0x56, 0x2A, 0x3E, 0x07, 0x20,
	0x15, 0x16, 0x26, 0x01, 0x20, 0x00, 0x05, 0x0C, 0x29, 0x2D, 0x4E, 0x27,
	0x0E, 0x1B, 0x2E, 0x05, 0x26, 0x5F, 0x03, 0x3C, 0x2C, 0x3F, 0x44, 0x2D,
	0x2F, 0x08, 0x2B, 0x21, 0x18, 0x2D, 0x29, 0x09, 0x06, 0x21, 0x0F, 0x24,
	0x05, 0x04, 0x00, 0x0F, 0x23, 0x00, 0x01, 0x3B, 0x2F, 0x38, 0x2B, 0x06,
	0x1B, 0x3E, 0x0C, 0x19, 0x40, 0x01, 0x01, 0x34, 0x2C, 0x0E, 0x13, 0x3F,
	0x30, 0x21, 0x2E, 0x0E, 0x54, 0x22, 0x08, 0x22, 0x29, 0x35, 0x25, 0x3A,
	0x58, 0x3A, 0x2A, 0x0E, 0x2A, 0x53, 0x25, 0x59, 0x06, 0x2D, 0x44, 0x24,
	0x29, 0x4A, 0x09, 0x02, 0x3B, 0x26, 0x36, 0x2F, 0x5C, 0x71, 0x58, 0x32,
	0x58, 0x27, 0x76, 0x3B, 0x07, 0x1D, 0x1A, 0x0A, 0x3E, 0x2D, 0x1A, 0x22,
	0x07, 0x02, 0x51, 0x2A, 0x1E, 0x10, 0x3E, 0x16, 0x1A, 0x39, 0x23, 0x26,
	0x26, 0x03, 0x03, 0x06, 0x23, 0x0E, 0x2A, 0x31, 0x7B, 0x39, 0x09, 0x05,
	0x2F, 0x16, 0x20, 0x26, 0x41, 0x3A, 0x1B, 0x07, 0x59, 0x09, 0x28, 0x77,
	0x28, 0x2D, 0x2A, 0x38, 0x29, 0x29, 0x30, 0x06, 0x22, 0x05, 0x21, 0x51,
	0x1F, 0x3E, 0x69, 0x05, 0x23, 0x24, 0x29, 0x77, 0x0B, 0x29, 0x2B, 0x25,
	0x11, 0x38, 0x30, 0x3D, 0x31, 0x03, 0x00, 0x06, 0x1E, 0x59, 0x1B, 0x07,
	0x18, 0x09, 0x23, 0x18, 0x2E, 0x05, 0x2D, 0x58, 0x0D, 0x35, 0x0A, 0x25,
	0x3A, 0x10, 0x35, 0x20, 0x41, 0x01, 0x13, 0x02, 0x34, 0x3F, 0x05, 0x0B,
	0x1D, 0x23, 0x39, 0x21, 0x21, 0x05, 0x50, 0x27, 0x0F, 0x03, 0x16, 0x0F,
	0x2C, 0x0D, 0x25, 0x27, 0x30, 0x04, 0x05, 0x0B, 0x2B, 0x2E, 0x23, 0x1F,
	0x11, 0x34, 0x30, 0x08, 0x31, 0x0B, 0x1B, 0x1B, 0x27, 0x3D, 0x11, 0x2F,
	0x0F, 0x2F, 0x3B, 0x1B, 0x1F, 0x30, 0x5D, 0x32, 0x01, 0x38, 0x2B, 0x29,
	0x2A, 0x13, 0x3D, 0x15, 0x26, 0x32, 0x30, 0x2B, 0x4A, 0x3C, 0x2A, 0x0F,
	0x3D, 0x02, 0x5A, 0x2F, 0x6D, 0x22, 0x14, 0x25, 0x39, 0x0F, 0x5D, 0x20,
	0x22, 0x0C, 0x17, 0x54, 0x22, 0x0D, 0x2E, 0x08, 0x59, 0x25, 0x22, 0x2A,
	0x33, 0x14, 0x23, 0x0D, 0x3A, 0x09, 0x58, 0x20, 0x28, 0x27, 0x13, 0x00,
	0x0A, 0x3F, 0x40, 0x0D, 0x2F, 0x53, 0x06, 0x05, 0x06, 0x3B, 0x34, 0x2C,
	0x2C, 0x23, 0x23, 0x0C, 0x2A, 0x32, 0x29, 0x05, 0x30, 0x0D, 0x32, 0x1B,
	0x2F, 0x22, 0x2B, 0x21, 0x18, 0x25, 0x1B, 0x02, 0x0D, 0x00, 0x25, 0x2F,
	0x2F, 0x13, 0x2C, 0x06, 0x18, 0x2F, 0x5F, 0x29, 0x01, 0x06, 0x2C, 0x12,
	0x0C, 0x19, 0x23, 0x3A, 0x28, 0x06, 0x07, 0x06, 0x37, 0x59, 0x3A, 0x0B,
	0x35, 0x58, 0x22, 0x2E, 0x25, 0x31, 0x23, 0x2A, 0x71, 0x3E, 0x53, 0x09,
	0x1D, 0x06, 0x04, 0x58, 0x19, 0x25, 0x21, 0x3D, 0x15, 0x01, 0x28, 0x0F,
	0x0F, 0x37, 0x23, 0x05, 0x07, 0x1C, 0x36, 0x2D, 0x01, 0x0E, 0x2A, 0x52,
	0x34, 0x13, 0x09, 0x08, 0x20, 0x06, 0x07, 0x28, 0x0B, 0x22, 0x3E, 0x00,
	0x25, 0x0A, 0x34, 0x2C, 0x3F, 0x72, 0x2B, 0x55, 0x2A, 0x11, 0x08, 0x2B,
	0x12, 0x3C, 0x24, 0x17, 0x24, 0x36, 0x3D, 0x26, 0x75, 0x0E, 0x15, 0x2F,
	0x59, 0x17, 0x24, 0x26, 0x21, 0x2A, 0x09, 0x2F, 0x0D, 0x07, 0x5E, 0x04,
	0x58, 0x51, 0x05, 0x22, 0x06, 0x39, 0x25, 0x29, 0x06, 0x0D, 0x00, 0x2C,
	0x27, 0x03, 0x75, 0x25, 0x26, 0x20, 0x0F, 0x01, 0x1F, 0x20, 0x37, 0x31,
	0x1B, 0x5B, 0x2E, 0x1B, 0x5F, 0x03, 0x09, 0x30, 0x23, 0x33, 0x74, 0x24,
	0x55, 0x2F, 0x2C, 0x3B, 0x3F, 0x1B, 0x0D, 0x38, 0x16, 0x09, 0x51, 0x2C,
	0x1D, 0x25, 0x2D, 0x54, 0x2C, 0x44, 0x03, 0x0F, 0x09, 0x28, 0x02, 0x13,
	0x27, 0x16, 0x2F, 0x5C, 0x7B, 0x05, 0x32, 0x3C, 0x29, 0x0D, 0x1F, 0x20,
	0x02, 0x00, 0x0B, 0x35, 0x22, 0x3A, 0x21, 0x05, 0x2A, 0x19, 0x0D, 0x38,
	0x16, 0x0F, 0x28, 0x56, 0x32, 0x06, 0x27, 0x24, 0x36, 0x21, 0x03, 0x14,
	0x54, 0x1B, 0x2E, 0x03, 0x21, 0x12, 0x0F, 0x27, 0x07, 0x22, 0x00, 0x2C,
	0x01, 0x12, 0x29, 0x53, 0x06, 0x29, 0x72, 0x0B, 0x38, 0x5C, 0x11, 0x2A,
	0x2F, 0x0C, 0x03, 0x29, 0x28, 0x22, 0x24, 0x0B, 0x1C, 0x2B, 0x01, 0x30,
	0x23, 0x3E, 0x74, 0x29, 0x34, 0x2F, 0x5E, 0x3B, 0x18, 0x06, 0x0B, 0x3E,
	0x00, 0x0F, 0x2B, 0x57, 0x09, 0x0B, 0x54, 0x52, 0x07, 0x39, 0x18, 0x2E,
	0x57, 0x2F, 0x52, 0x28, 0x28, 0x12, 0x34, 0x3D, 0x07, 0x27, 0x33, 0x5A,
	0x19, 0x03, 0x3C, 0x02, 0x2D, 0x1A, 0x04, 0x3F, 0x37, 0x41, 0x05, 0x30,
	0x2D, 0x13, 0x45, 0x58, 0x6D, 0x55, 0x12, 0x5C, 0x3A, 0x2D, 0x5D, 0x34,
	0x38, 0x5D, 0x0F, 0x25, 0x20, 0x0F, 0x2D, 0x04, 0x1D, 0x36, 0x18, 0x31,
	0x1B, 0x1B, 0x0C, 0x18, 0x44, 0x13, 0x14, 0x18, 0x1D, 0x2E, 0x38, 0x3B,
	0x3B, 0x1D, 0x00, 0x77, 0x1E, 0x10, 0x3A, 0x18, 0x70, 0x3D, 0x14, 0x37,
	0x52, 0x77, 0x1F, 0x00, 0x5E, 0x09, 0x6D, 0x18, 0x51, 0x28, 0x02, 0x16,
	0x06, 0x06, 0x3E, 0x1C, 0x34, 0x3E, 0x06, 0x0A, 0x01, 0x0B, 0x3F, 0x14,
	0x03, 0x19, 0x2D, 0x19, 0x51, 0x3F, 0x11, 0x14, 0x01, 0x27, 0x0A, 0x52,
	0x10, 0x18, 0x3B, 0x38, 0x53, 0x7B, 0x3F, 0x0D, 0x20, 0x26, 0x23, 0x3E,
	0x07, 0x2D, 0x3E, 0x26, 0x14, 0x28, 0x3C, 0x5D, 0x05, 0x04, 0x03, 0x5F,
	0x20, 0x01, 0x5C, 0x52, 0x20, 0x3F, 0x76, 0x3A, 0x32, 0x3B, 0x1B, 0x33,
	0x5C, 0x07, 0x05, 0x58, 0x03, 0x54, 0x19, 0x14, 0x20, 0x06, 0x58, 0x3B,
	0x3D, 0x0E, 0x00, 0x1A, 0x51, 0x29, 0x1A, 0x32, 0x03, 0x57, 0x1F, 0x08,
	0x7A, 0x08, 0x13, 0x37, 0x06, 0x29, 0x06, 0x31, 0x3A, 0x32, 0x37, 0x1A,
	0x26, 0x0F, 0x00, 0x2A, 0x39, 0x33, 0x0B, 0x04, 0x2E, 0x36, 0x2B, 0x02,
	0x3F, 0x00, 0x1B, 0x38, 0x5D, 0x5C, 0x17, 0x25, 0x36, 0x57, 0x07, 0x23,
	0x5E, 0x03, 0x3C, 0x18, 0x0B, 0x1C, 0x31, 0x06, 0x58, 0x07, 0x01, 0x39,
	0x22, 0x29, 0x08, 0x07, 0x05, 0x3C, 0x20, 0x32, 0x5E, 0x19, 0x20, 0x53,
	0x13, 0x00, 0x12, 0x20, 0x0A, 0x10, 0x21, 0x2F, 0x2B, 0x09, 0x03, 0x3F,
	0x0C, 0x00, 0x1F, 0x06, 0x54, 0x2E, 0x05, 0x5B, 0x76, 0x3C, 0x18, 0x2F,
	0x25, 0x27, 0x07, 0x55, 0x0C, 0x00, 0x35, 0x0F, 0x2D, 0x2B, 0x08, 0x38,
	0x1F, 0x13, 0x27, 0x1F, 0x11, 0x26, 0x27, 0x5D, 0x07, 0x11, 0x55, 0x13,
	0x5E, 0x07, 0x0A, 0x01, 0x26, 0x03, 0x06, 0x32, 0x22, 0x18, 0x25, 0x06,
	0x29, 0x3C, 0x13, 0x56, 0x0E, 0x32, 0x2A, 0x57, 0x2B, 0x1F, 0x73, 0x3F,
	0x03, 0x38, 0x1C, 0x71, 0x2E, 0x2C, 0x29, 0x12, 0x24, 0x3A, 0x2A, 0x38,
	0x5C, 0x1B, 0x1D, 0x59, 0x39, 0x09, 0x3B, 0x54, 0x29, 0x2B, 0x02, 0x08,
	0x5D, 0x50, 0x3C, 0x2F, 0x2F, 0x1A, 0x38, 0x17, 0x11, 0x3A, 0x2B, 0x26,
	0x5C, 0x18, 0x28, 0x1B, 0x06, 0x2C, 0x5E, 0x24, 0x22, 0x50, 0x24, 0x23,
	0x2D, 0x05, 0x52, 0x3F, 0x20, 0x36, 0x39, 0x0E, 0x3B, 0x5D, 0x31, 0x0B,
	0x38, 0x36, 0x5E, 0x06, 0x5A, 0x26, 0x1D, 0x03, 0x24, 0x34, 0x12, 0x0A,
	0x1D, 0x2C, 0x0D, 0x0A, 0x02, 0x00, 0x10, 0x38, 0x0E, 0x28, 0x2C, 0x33,
	0x3A, 0x0A, 0x34, 0x3C, 0x09, 0x22, 0x2A, 0x1C, 0x12, 0x20, 0x09, 0x57,
	0x29, 0x1E, 0x33, 0x5A, 0x51, 0x34, 0x1B, 0x7A, 0x06, 0x34, 0x06, 0x5A,
	0x01, 0x08, 0x53, 0x29, 0x08, 0x0E, 0x1C, 0x14, 0x20, 0x0A, 0x11, 0x20,
	0x4A, 0x0B, 0x0C, 0x23, 0x09, 0x2D, 0x34, 0x25, 0x33, 0x26, 0x03, 0x58,
	0x32, 0x6D, 0x19, 0x03, 0x59, 0x03, 0x31, 0x29, 0x34, 0x01, 0x3B, 0x77,
	0x3C, 0x0C, 0x29, 0x18, 0x25, 0x58, 0x16, 0x24, 0x3E, 0x74, 0x3F, 0x02,
	0x25, 0x1A, 0x05, 0x06, 0x06, 0x36, 0x3F, 0x31, 0x22, 0x07, 0x04, 0x1A,
	0x29, 0x3B, 0x0E, 0x3D, 0x38, 0x29, 0x2F, 0x36, 0x09, 0x1B, 0x74, 0x5A,
	0x59, 0x3F, 0x2E, 0x06, 0x1A, 0x0F, 0x5B, 0x00, 0x12, 0x35, 0x0D, 0x0B,
	0x1A, 0x17, 0x5A, 0x3B, 0x38, 0x04, 0x14, 0x2B, 0x11, 0x0F, 0x12, 0x7B,
	0x27, 0x4E, 0x02, 0x0F, 0x27, 0x0E, 0x4A, 0x0B, 0x1B, 0x2C, 0x1D, 0x58,
	0x37, 0x2C, 0x70, 0x47, 0x37, 0x1F, 0x38, 0x2F, 0x2E, 0x25, 0x19, 0x03,
	0x33, 0x16, 0x58, 0x1A, 0x0F, 0x23, 0x38, 0x15, 0x1E, 0x18, 0x77, 0x34,
	0x08, 0x58, 0x3A, 0x29, 0x36, 0x28, 0x36, 0x08, 0x2A, 0x19, 0x39, 0x38,
	0x09, 0x23, 0x05, 0x11, 0x26, 0x22, 0x73, 0x5C, 0x0E, 0x38, 0x5D, 0x0C,
	0x39, 0x39, 0x38, 0x27, 0x2E, 0x21, 0x10, 0x01, 0x09, 0x07, 0x08, 0x15,
	0x3E, 0x1A, 0x1A, 0x38, 0x36, 0x5F, 0x07, 0x38, 0x09, 0x0F, 0x36, 0x3D,
	0x35, 0x5B, 0x06, 0x0F, 0x0E, 0x01, 0x22, 0x15, 0x34, 0x2E, 0x10, 0x35,
	0x28, 0x5C, 0x5C, 0x0C, 0x1D, 0x56, 0x2D, 0x5E, 0x23, 0x38, 0x52, 0x3B,
	0x0F, 0x08, 0x0B, 0x26, 0x0F, 0x1B, 0x2B, 0x0B, 0x0B, 0x09, 0x11, 0x34,
	0x5D, 0x11, 0x2C, 0x06, 0x16, 0x0A, 0x57, 0x3A, 0x5A, 0x3A, 0x5C, 0x14,
	0x37, 0x11, 0x11, 0x1E, 0x0B, 0x22, 0x3A, 0x24, 0x16, 0x00, 0x1C, 0x5C,
	0x31, 0x0E, 0x38, 0x58, 0x13, 0x37, 0x5C, 0x0C, 0x04, 0x3C, 0x29, 0x5F,
	0x15, 0x27, 0x5E, 0x3A, 0x20, 0x39, 0x29, 0x25, 0x33, 0x1A, 0x31, 0x5A,
	0x0A, 0x27, 0x58, 0x30, 0x22, 0x09, 0x2A, 0x58, 0x51, 0x37, 0x38, 0x0E,
	0x21, 0x06, 0x5E, 0x32, 0x04, 0x22, 0x34, 0x3C, 0x2C, 0x2D, 0x0A, 0x03,
	0x02, 0x1D, 0x04, 0x1D, 0x33, 0x25, 0x2D, 0x71, 0x14, 0x0F, 0x2F, 0x31,
	0x17, 0x2E, 0x59, 0x1B, 0x18, 0x70, 0x2E, 0x55, 0x3E, 0x2C, 0x13, 0x25,
	0x0C, 0x09, 0x5A, 0x03, 0x5C, 0x16, 0x2F, 0x5B, 0x7B, 0x39, 0x26, 0x14,
	0x23, 0x33, 0x0B, 0x11, 0x00, 0x1A, 0x70, 0x38, 0x58, 0x5E, 0x07, 0x2E,
	0x36, 0x28, 0x57, 0x3D, 0x7A, 0x1A, 0x2B, 0x1F, 0x1C, 0x34, 0x1B, 0x2A,
	0x0C, 0x2D, 0x0A, 0x1F, 0x28, 0x58, 0x3C, 0x70, 0x16, 0x53, 0x00, 0x3F,
	0x16, 0x0D, 0x13, 0x0C, 0x5C, 0x0C, 0x29, 0x20, 0x0B, 0x39, 0x13, 0x09,
	0x2B, 0x1C, 0x18, 0x37, 0x23, 0x24, 0x3A, 0x0A, 0x16, 0x16, 0x11, 0x27,
	0x1F, 0x2A, 0x5D, 0x53, 0x09, 0x2F, 0x10, 0x20, 0x53, 0x2B, 0x53, 0x70,
	0x25, 0x00, 0x0F, 0x19, 0x05, 0x43, 0x24, 0x20, 0x22, 0x35, 0x5C, 0x0A,
	0x45, 0x04, 0x08, 0x5A, 0x11, 0x0C, 0x1B, 0x2E, 0x5E, 0x0F, 0x3A, 0x5E,
	0x21, 0x28, 0x4E, 0x39, 0x3D, 0x0C, 0x0F, 0x29, 0x00, 0x5A, 0x16, 0x5D,
	0x35, 0x21, 0x29, 0x35, 0x1A, 0x52, 0x04, 0x2F, 0x74, 0x04, 0x02, 0x5F,
	0x5D, 0x26, 0x2F, 0x02, 0x05, 0x3C, 0x33, 0x23, 0x03, 0x3A, 0x1F, 0x75,
	0x24, 0x27, 0x22, 0x1E, 0x27, 0x5A, 0x03, 0x0F, 0x12, 0x06, 0x3F, 0x09,
	0x23, 0x3C, 0x04, 0x21, 0x59, 0x2B, 0x07, 0x26, 0x1A, 0x0A, 0x58, 0x00,
	0x36, 0x07, 0x30, 0x22, 0x3C, 0x09, 0x0D, 0x07, 0x04, 0x5A, 0x12, 0x1D,
	0x29, 0x17, 0x5A, 0x73, 0x39, 0x02, 0x1D, 0x2E, 0x26, 0x0E, 0x39, 0x29,
	0x03, 0x08, 0x58, 0x36, 0x5E, 0x52, 0x76, 0x29, 0x2C, 0x3E, 0x19, 0x08,
	0x5E, 0x14, 0x29, 0x3A, 0x04, 0x01, 0x0B, 0x27, 0x1B, 0x70, 0x58, 0x00,
	0x2D, 0x32, 0x69, 0x5B, 0x00, 0x01, 0x01, 0x09, 0x02, 0x35, 0x36, 0x28,
	0x28, 0x02, 0x39, 0x3C, 0x28, 0x0C, 0x06, 0x09, 0x1E, 0x24, 0x04, 0x3E,
	0x57, 0x25, 0x01, 0x10, 0x08, 0x34, 0x28, 0x05, 0x06, 0x0A, 0x15, 0x24,
	0x05, 0x16, 0x38, 0x00, 0x2A, 0x05, 0x12, 0x3D, 0x2C, 0x2B, 0x1D, 0x2D,
	0x1D, 0x2F, 0x29, 0x2E, 0x05, 0x27, 0x27, 0x36, 0x11, 0x11, 0x08, 0x18,
	0x41, 0x5E, 0x30, 0x1D, 0x06, 0x3A, 0x58, 0x1B, 0x14, 0x55, 0x5F, 0x19,
	0x23, 0x3F, 0x58, 0x0A, 0x1A, 0x6D, 0x3C, 0x12, 0x21, 0x1A, 0x37, 0x1C,
	0x39, 0x57, 0x0D, 0x15, 0x1C, 0x16, 0x17, 0x5A, 0x73, 0x2D, 0x51, 0x24,
	0x38, 0x7A, 0x38, 0x14, 0x2F, 0x3F, 0x15, 0x23, 0x13, 0x57, 0x02, 0x1A,
	0x1F, 0x19, 0x02, 0x0D, 0x09, 0x1A, 0x14, 0x18, 0x19, 0x2F, 0x23, 0x50,
	0x57, 0x33, 0x04, 0x5E, 0x52, 0x3D, 0x02, 0x12, 0x47, 0x35, 0x36, 0x31,
	0x2B, 0x09, 0x0E, 0x37, 0x27, 0x3A, 0x2E, 0x1B, 0x3A, 0x00, 0x2A, 0x38,
	0x12, 0x1E, 0x05, 0x70, 0x03, 0x53, 0x59, 0x25, 0x20, 0x0E, 0x36, 0x5C,
	0x08, 0x76, 0x1A, 0x18, 0x1B, 0x2D, 0x18, 0x0E, 0x17, 0x58, 0x58, 0x36,
	0x34, 0x27, 0x29, 0x33, 0x24, 0x07, 0x52, 0x02, 0x5B, 0x36, 0x22, 0x20,
	0x0B, 0x0C, 0x2C, 0x3D, 0x56, 0x5A, 0x20, 0x18, 0x54, 0x15, 0x0A, 0x3E,
	0x26, 0x1B, 0x3B, 0x0F, 0x12, 0x03, 0x28, 0x00, 0x20, 0x1B, 0x37, 0x3A,
	0x02, 0x3D, 0x59, 0x77, 0x34, 0x26, 0x5E, 0x59, 0x76, 0x34, 0x2F, 0x04,
	0x26, 0x08, 0x1B, 0x03, 0x08, 0x5C, 0x1A, 0x21, 0x15, 0x0D, 0x11, 0x2C,
	0x0D, 0x14, 0x38, 0x19, 0x2F, 0x0B, 0x04, 0x0F, 0x5D, 0x2D, 0x0D, 0x00,
	0x3A, 0x1F, 0x08, 0x29, 0x0B, 0x39, 0x2F, 0x31, 0x1E, 0x30, 0x57, 0x01,
	0x30, 0x16, 0x57, 0x02, 0x2F, 0x11, 0x34, 0x20, 0x1D, 0x11, 0x0D, 0x3B,
	0x17, 0x06, 0x13, 0x73, 0x5D, 0x35, 0x1C, 0x29, 0x71, 0x2F, 0x50, 0x0F,
	0x26, 0x1A, 0x0A, 0x03, 0x57, 0x2A, 0x36, 0x59, 0x17, 0x58, 0x07, 0x04,
	0x36, 0x56, 0x37, 0x20, 0x15, 0x43, 0x59, 0x3A, 0x59, 0x20, 0x58, 0x36,
	0x21, 0x0E, 0x72, 0x34, 0x55, 0x1A, 0x0A, 0x2F, 0x07, 0x50, 0x0F, 0x2F,
	0x38, 0x3D, 0x00, 0x0F, 0x05, 0x13, 0x1B, 0x0E, 0x00, 0x3C, 0x01, 0x01,
	0x58, 0x5B, 0x38, 0x33, 0x06, 0x27, 0x0B, 0x09, 0x1A, 0x0D, 0x13, 0x05,
	0x59, 0x37, 0x0E, 0x15, 0x1F, 0x18, 0x33, 0x01, 0x2F, 0x3E, 0x40, 0x12,
	0x22, 0x00, 0x16, 0x0A, 0x13, 0x02, 0x15, 0x05, 0x2C, 0x35, 0x5F, 0x34,
	0x1C, 0x31, 0x07, 0x2B, 0x0A, 0x1C, 0x20, 0x76, 0x05, 0x50, 0x37, 0x0A,
	0x3B, 0x2E, 0x59, 0x5A, 0x3B, 0x27, 0x21, 0x10, 0x3A, 0x1F, 0x08, 0x23,
	0x20, 0x57, 0x5B, 0x71, 0x5C, 0x34, 0x2A, 0x3C, 0x28, 0x0D, 0x10, 0x5A,
	0x28, 0x21, 0x2F, 0x11, 0x20, 0x3D, 0x0C, 0x09, 0x0B, 0x02, 0x1E, 0x70,
	0x22, 0x37, 0x2A, 0x02, 0x15, 0x16, 0x31, 0x59, 0x09, 0x25, 0x1B, 0x2A,
	0x29, 0x24, 0x38, 0x3C, 0x0E, 0x27, 0x3F, 0x00, 0x5C, 0x30, 0x16, 0x24,
	0x1B, 0x5F, 0x20, 0x1E, 0x0C, 0x69, 0x1F, 0x38, 0x5D, 0x26, 0x24, 0x0B,
	0x33, 0x3F, 0x09, 0x34, 0x21, 0x4E, 0x07, 0x2C, 0x13, 0x36, 0x52, 0x03,
	0x26, 0x2F, 0x16, 0x26, 0x01, 0x2A, 0x0D, 0x28, 0x03, 0x09, 0x1C, 0x0D,
	0x36, 0x29, 0x2F, 0x04, 0x25, 0x47, 0x2C, 0x37, 0x11, 0x05, 0x3A, 0x16,
	0x28, 0x32, 0x12, 0x0E, 0x26, 0x2D, 0x13, 0x28, 0x54, 0x23, 0x0F, 0x2F,
	0x1A, 0x14, 0x0B, 0x3B, 0x09, 0x3B, 0x2A, 0x25, 0x26, 0x04, 0x0D, 0x08,
	0x26, 0x0B, 0x11, 0x04, 0x58, 0x24, 0x2F, 0x2C, 0x32, 0x3D, 0x1B, 0x21,
	0x32, 0x0E, 0x2F, 0x30, 0x19, 0x33, 0x72, 0x21, 0x0F, 0x03, 0x0D, 0x35,
	0x21, 0x38, 0x20, 0x1A, 0x0E, 0x3B, 0x37, 0x01, 0x1C, 0x33, 0x2D, 0x37,
	0x09, 0x11, 0x72, 0x35, 0x25, 0x29, 0x2E, 0x35, 0x0B, 0x02, 0x26, 0x03,
	0x06, 0x29, 0x54, 0x04, 0x08, 0x03, 0x01, 0x25, 0x58, 0x13, 0x25, 0x54,
	0x16, 0x1B, 0x2A, 0x73, 0x2E, 0x11, 0x56, 0x12, 0x69, 0x25, 0x0D, 0x2C,
	0x2F, 0x18, 0x58, 0x2C, 0x14, 0x39, 0x2C, 0x1F, 0x1B, 0x29, 0x2A, 0x25,
	0x0B, 0x16, 0x23, 0x31, 0x16, 0x2B, 0x27, 0x19, 0x2A, 0x2D, 0x23, 0x54,
	0x2A, 0x29, 0x1B, 0x16, 0x04, 0x27, 0x27, 0x00, 0x0D, 0x16, 0x19, 0x40,
	0x18, 0x3C, 0x20, 0x22, 0x0C, 0x38, 0x1C, 0x0C, 0x3A, 0x27, 0x72, 0x1B,
	0x00, 0x23, 0x40, 0x25, 0x2E, 0x55, 0x3E, 0x52, 0x05, 0x39, 0x19, 0x07,
	0x08, 0x03, 0x1D, 0x25, 0x1D, 0x13, 0x2E, 0x0F, 0x16, 0x0B, 0x2A, 0x2A,
	0x2E, 0x12, 0x1D, 0x31, 0x24, 0x21, 0x0B, 0x09, 0x29, 0x35, 0x0E, 0x37,
	0x14, 0x2C, 0x1A, 0x35, 0x08, 0x2B, 0x2D, 0x0E, 0x2E, 0x13, 0x1D, 0x13,
	0x05, 0x2B, 0x1B, 0x21, 0x09, 0x18, 0x0F, 0x25, 0x03, 0x0D, 0x70, 0x04,
	0x25, 0x2B, 0x5E, 0x2B, 0x0F, 0x23, 0x58, 0x2F, 0x3A, 0x3D, 0x1B, 0x1B,
	0x32, 0x24, 0x2D, 0x24, 0x09, 0x40, 0x17, 0x21, 0x31, 0x03, 0x09, 0x35,
	0x29, 0x55, 0x23, 0x0A, 0x30, 0x3B, 0x35, 0x37, 0x0C, 0x0F, 0x24, 0x36,
	0x2A, 0x2F, 0x2D, 0x14, 0x26, 0x23, 0x13, 0x25, 0x2F, 0x0E, 0x21, 0x3F,
	0x05, 0x26, 0x1B, 0x26, 0x5F, 0x03, 0x03, 0x26, 0x1A, 0x11, 0x01, 0x58,
	0x0B, 0x56, 0x2D, 0x28, 0x28, 0x27, 0x5B, 0x00, 0x7A, 0x2E, 0x00, 0x2A,
	0x05, 0x3A, 0x0B, 0x51, 0x0C, 0x26, 0x70, 0x39, 0x0D, 0x5E, 0x2E, 0x0A,
	0x2E, 0x0B, 0x5E, 0x32, 0x06, 0x2B, 0x30, 0x19, 0x0C, 0x31, 0x2A, 0x0E,
	0x2C, 0x1B, 0x0F, 0x35, 0x29, 0x23, 0x19, 0x25, 0x23, 0x20, 0x34, 0x11,
	0x05, 0x3A, 0x1B, 0x25, 0x32, 0x00, 0x2B, 0x25, 0x1E, 0x13, 0x2A, 0x54,
	0x1B, 0x1B, 0x2A, 0x2C, 0x2E, 0x13, 0x3B, 0x18, 0x2F, 0x24, 0x28, 0x14,
	0x59, 0x0B, 0x14, 0x23, 0x3D, 0x1C, 0x18, 0x18, 0x26, 0x0B, 0x11, 0x00,
	0x35, 0x22, 0x3D, 0x2F, 0x07, 0x0B, 0x00, 0x26, 0x26, 0x38, 0x05, 0x23,
	0x19, 0x39, 0x29, 0x21, 0x2D, 0x03, 0x22, 0x35, 0x02, 0x59, 0x2B, 0x38,
	0x00, 0x02, 0x02, 0x16, 0x0E, 0x0B, 0x38, 0x23, 0x56, 0x1C, 0x38, 0x09,
	0x38, 0x18, 0x2A, 0x32, 0x0B, 0x19, 0x56, 0x32, 0x10, 0x26, 0x38, 0x17,
	0x5A, 0x05, 0x3C, 0x30, 0x06, 0x2E, 0x07, 0x09, 0x06, 0x5F, 0x32, 0x0F,
	0x54, 0x09, 0x02, 0x5B, 0x18, 0x18, 0x22, 0x20, 0x3A, 0x1A, 0x54, 0x26,
	0x3F, 0x13, 0x25, 0x0F, 0x18, 0x29, 0x2A, 0x01, 0x0B, 0x19, 0x27, 0x2C,
	0x2A, 0x16, 0x26, 0x37, 0x11, 0x27, 0x2D, 0x34, 0x2C, 0x06, 0x21, 0x16,
	0x14, 0x27, 0x01, 0x00, 0x3A, 0x30, 0x17, 0x1E, 0x1B, 0x5F, 0x20, 0x0C,
	0x0C, 0x74, 0x39, 0x2C, 0x00, 0x06, 0x06, 0x1B, 0x28, 0x01, 0x24, 0x71,
	0x2B, 0x29, 0x14, 0x26, 0x76, 0x2E, 0x12, 0x29, 0x1D, 0x38, 0x2B, 0x0E,
	0x5E, 0x3E, 0x23, 0x2B, 0x4A, 0x09, 0x12, 0x23, 0x21, 0x26, 0x04, 0x24,
	0x2D, 0x28, 0x36, 0x2A, 0x05, 0x10, 0x00, 0x51, 0x37, 0x0F, 0x01, 0x0A,
	0x16, 0x3A, 0x2A, 0x05, 0x25, 0x58, 0x1A, 0x1C, 0x69, 0x54, 0x02, 0x09,
	0x1B, 0x24, 0x5F, 0x07, 0x5A, 0x5C, 0x2D, 0x21, 0x07, 0x5A, 0x44, 0x30,
	0x38, 0x2D, 0x5D, 0x53, 0x0A, 0x18, 0x05, 0x02, 0x40, 0x24, 0x54, 0x04,
	0x5F, 0x59, 0x2C, 0x54, 0x31, 0x0F, 0x5F, 0x38, 0x43, 0x07, 0x3C, 0x44,
	0x70, 0x0E, 0x06, 0x0B, 0x1A, 0x69, 0x58, 0x15, 0x02, 0x04, 0x23, 0x01,
	0x08, 0x57, 0x26, 0x01, 0x03, 0x54, 0x22, 0x2D, 0x76, 0x0A, 0x06, 0x34,
	0x22, 0x0C, 0x0A, 0x38, 0x5C, 0x2F, 0x00, 0x14, 0x0B, 0x2A, 0x3A, 0x73,
	0x06, 0x07, 0x38, 0x29, 0x21, 0x18, 0x0C, 0x36, 0x18, 0x36, 0x3C, 0x30,
	0x0A, 0x24, 0x11, 0x09, 0x0D, 0x24, 0x19, 0x0D, 0x0A, 0x25, 0x09, 0x09,
	0x20, 0x39, 0x31, 0x1B, 0x1A, 0x18, 0x25, 0x12, 0x1C, 0x53, 0x13, 0x07,
	0x08, 0x26, 0x0C, 0x13, 0x19, 0x00, 0x08, 0x03, 0x04, 0x47, 0x02, 0x57,
	0x2E, 0x36, 0x3C, 0x0E, 0x17, 0x2D, 0x2C, 0x04, 0x4A, 0x24, 0x00, 0x26,
	0x2B, 0x38, 0x0D, 0x5A, 0x1A, 0x22, 0x27, 0x28, 0x5A, 0x2E, 0x58, 0x55,
	0x25, 0x06, 0x24, 0x5E, 0x07, 0x25, 0x27, 0x11, 0x35, 0x17, 0x5E, 0x3F,
	0x17, 0x1B, 0x00, 0x26, 0x04, 0x72, 0x0F, 0x2C, 0x27, 0x5B, 0x2B, 0x39,
	0x08, 0x2C, 0x2D, 0x74, 0x26, 0x05, 0x57, 0x27, 0x11, 0x58, 0x51, 0x3C,
	0x1B, 0x74, 0x08, 0x25, 0x0F, 0x07, 0x7A, 0x35, 0x33, 0x1E, 0x02, 0x14,
	0x24, 0x2B, 0x5C, 0x0A, 0x2E, 0x2E, 0x06, 0x04, 0x02, 0x6D, 0x3B, 0x2F,
	0x37, 0x3E, 0x0C, 0x07, 0x0F, 0x45, 0x31, 0x05, 0x3E, 0x0E, 0x3D, 0x23,
	0x0D, 0x28, 0x0E, 0x04, 0x58, 0x25, 0x5F, 0x53, 0x2C, 0x02, 0x0C, 0x07,
	0x22, 0x00, 0x1F, 0x08, 0x35, 0x10, 0x00, 0x32, 0x12, 0x3F, 0x50, 0x3C,
	0x06, 0x2A, 0x0B, 0x35, 0x02, 0x08, 0x11, 0x54, 0x14, 0x37, 0x59, 0x74,
	0x29, 0x24, 0x01, 0x0D, 0x03, 0x39, 0x02, 0x57, 0x28, 0x21, 0x54, 0x34,
	0x1F, 0x3F, 0x2A, 0x22, 0x36, 0x3C, 0x2C, 0x2E, 0x29, 0x11, 0x59, 0x2F,
	0x07, 0x1D, 0x39, 0x17, 0x5A, 0x0C, 0x22, 0x06, 0x3A, 0x1C, 0x0B, 0x3E,
	0x31, 0x25, 0x18, 0x69, 0x35, 0x22, 0x45, 0x00, 0x71, 0x5D, 0x38, 0x29,
	0x2A, 0x76, 0x0F, 0x35, 0x1B, 0x2C, 0x16, 0x58, 0x39, 0x08, 0x0E, 0x13,
	0x3A, 0x26, 0x28, 0x3C, 0x37, 0x00, 0x32, 0x0D, 0x01, 0x05, 0x3B, 0x24,
	0x24, 0x0C, 0x09, 0x0A, 0x24, 0x05, 0x1D, 0x75, 0x28, 0x04, 0x36, 0x3A,
	0x31, 0x00, 0x05, 0x07, 0x3C, 0x30, 0x1C, 0x34, 0x5B, 0x0C, 0x23, 0x5C,
	0x09, 0x29, 0x32, 0x01, 0x14, 0x02, 0x23, 0x32, 0x1B, 0x06, 0x17, 0x06,
	0x03, 0x14, 0x47, 0x4A, 0x02, 0x0C, 0x18, 0x2D, 0x0E, 0x0F, 0x3B, 0x2B,
	0x1F, 0x02, 0x37, 0x1E, 0x03, 0x1E, 0x59, 0x41, 0x33, 0x2E, 0x23, 0x2E,
	0x1B, 0x40, 0x29, 0x06, 0x4E, 0x01, 0x05, 0x10, 0x47, 0x2D, 0x5F, 0x5F,
	0x36, 0x26, 0x4E, 0x19, 0x2D, 0x33, 0x09, 0x28, 0x5E, 0x5D, 0x00, 0x25,
	0x56, 0x1F, 0x00, 0x32, 0x5A, 0x00, 0x02, 0x21, 0x1B, 0x02, 0x05, 0x1E,
	0x3C, 0x32, 0x20, 0x0F, 0x3B, 0x22, 0x2B, 0x2D, 0x34, 0x2D, 0x3E, 0x21,
	0x07, 0x56, 0x1F, 0x05, 0x08, 0x07, 0x12, 0x17, 0x1B, 0x0B, 0x1D, 0x00,
	0x1C, 0x00, 0x24, 0x3F, 0x29, 0x25, 0x5B, 0x23, 0x07, 0x23, 0x01, 0x27,
	0x2E, 0x04, 0x10, 0x16, 0x06, 0x09, 0x2D, 0x2C, 0x25, 0x38, 0x2B, 0x5B,
	0x16, 0x5F, 0x3C, 0x29, 0x2A, 0x02, 0x5D, 0x20, 0x71, 0x05, 0x54, 0x03,
	0x0A, 0x25, 0x22, 0x3B, 0x1D, 0x11, 0x2B, 0x59, 0x03, 0x5C, 0x12, 0x33,
	0x0F, 0x03, 0x59, 0x2A, 0x69, 0x01, 0x26, 0x5C, 0x21, 0x37, 0x23, 0x33,
	0x18, 0x52, 0x09, 0x3E, 0x12, 0x25, 0x02, 0x72, 0x3E, 0x31, 0x16, 0x5E,
	0x18, 0x3A, 0x02, 0x05, 0x04, 0x0B, 0x47, 0x20, 0x5C, 0x52, 0x71, 0x2E,
	0x2D, 0x26, 0x06, 0x15, 0x1D, 0x25, 0x0B, 0x09, 0x18, 0x38, 0x2D, 0x1A,
	0x03, 0x38, 0x01, 0x57, 0x0B, 0x3E, 0x29, 0x04, 0x52, 0x39, 0x0C, 0x2D,
	0x24, 0x34, 0x5A, 0x5E, 0x16, 0x1F, 0x00, 0x03, 0x39, 0x01, 0x39, 0x2B,
	0x01, 0x1A, 0x13, 0x26, 0x14, 0x22, 0x03, 0x37, 0x3B, 0x03, 0x24, 0x1A,
	0x06, 0x07, 0x04, 0x1E, 0x52, 0x0E, 0x2B, 0x2C, 0x24, 0x26, 0x17, 0x04,
	0x51, 0x2C, 0x40, 0x09, 0x23, 0x07, 0x45, 0x04, 0x26, 0x27, 0x0C, 0x00,
	0x5C, 0x08, 0x34, 0x3B, 0x17, 0x33, 0x25, 0x0A, 0x39, 0x24, 0x20, 0x10,
	0x3E, 0x25, 0x0A, 0x3C, 0x30, 0x23, 0x34, 0x25, 0x3B, 0x20, 0x54, 0x57,
	0x2D, 0x58, 0x05, 0x02, 0x37, 0x1C, 0x2C, 0x3B, 0x20, 0x24, 0x2A, 0x11,
	0x01, 0x23, 0x00, 0x19, 0x58, 0x21, 0x1B, 0x2D, 0x1D, 0x0D, 0x2B, 0x26,
	0x28, 0x29, 0x28, 0x07, 0x09, 0x2F, 0x03, 0x2E, 0x06, 0x25, 0x0D, 0x18,
	0x38, 0x2E, 0x14, 0x10, 0x21, 0x23, 0x2D, 0x1D, 0x38, 0x5C, 0x20, 0x18,
	0x59, 0x0E, 0x0B, 0x40, 0x72, 0x1A, 0x15, 0x5E, 0x18, 0x7A, 0x29, 0x2A,
	0x07, 0x20, 0x03, 0x39, 0x4A, 0x59, 0x0C, 0x18, 0x19, 0x00, 0x0C, 0x27,
	0x05, 0x14, 0x02, 0x17, 0x1C, 0x07, 0x08, 0x0A, 0x5B, 0x32, 0x27, 0x5A,
	0x0A, 0x05, 0x27, 0x0E, 0x3D, 0x00, 0x09, 0x07, 0x38, 0x3F, 0x39, 0x29,
	0x2F, 0x0A, 0x0E, 0x29, 0x2D, 0x11, 0x1B, 0x0B, 0x54, 0x2B, 0x5A, 0x77,
	0x26, 0x57, 0x38, 0x2C, 0x0F, 0x1B, 0x15, 0x2B, 0x04, 0x07, 0x2E, 0x0C,
	0x2A, 0x5C, 0x21, 0x3B, 0x14, 0x3E, 0x20, 0x2C, 0x0A, 0x27, 0x23, 0x38,
	0x7A, 0x34, 0x17, 0x25, 0x02, 0x21, 0x23, 0x13, 0x57, 0x32, 0x31, 0x2A,
	0x0D, 0x29, 0x53, 0x74, 0x5F, 0x39, 0x41, 0x02, 0x3A, 0x3B, 0x0A, 0x2D,
	0x59, 0x26, 0x1A, 0x27, 0x1F, 0x21, 0x38, 0x15, 0x27, 0x5E, 0x08, 0x0C,
	0x1E, 0x00, 0x0F, 0x20, 0x20, 0x00, 0x25, 0x45, 0x1A, 0x14, 0x2B, 0x19,
	0x3A, 0x24, 0x37, 0x28, 0x34, 0x1A, 0x52, 0x2F, 0x5B, 0x55, 0x08, 0x01,
	0x32, 0x58, 0x34, 0x2D, 0x26, 0x32, 0x27, 0x0A, 0x07, 0x3C, 0x77, 0x36,
	0x51, 0x2A, 0x07, 0x16, 0x1B, 0x19, 0x20, 0x01, 0x3A, 0x09, 0x55, 0x24,
	0x3E, 0x15, 0x02, 0x28, 0x3C, 0x3E, 0x72, 0x0B, 0x27, 0x09, 0x44, 0x05,
	0x16, 0x0E, 0x1B, 0x07, 0x0D, 0x43, 0x11, 0x09, 0x25, 0x24, 0x1C, 0x0D,
	0x37, 0x2E, 0x0A, 0x3A, 0x51, 0x06, 0x03, 0x72, 0x29, 0x36, 0x2D, 0x18,
	0x11, 0x0D, 0x11, 0x5C, 0x13, 0x0B, 0x18, 0x04, 0x03, 0x38, 0x0B, 0x00,
	0x2B, 0x09, 0x1D, 0x0C, 0x3A, 0x20, 0x1B, 0x3C, 0x04, 0x3E, 0x59, 0x5D,
	0x3D, 0x21, 0x04, 0x13, 0x20, 0x19, 0x70, 0x3C, 0x39, 0x37, 0x3F, 0x13,
	0x3E, 0x11, 0x2D, 0x3F, 0x17, 0x58, 0x05, 0x17, 0x39, 0x33, 0x20, 0x25,
	0x19, 0x20, 0x14, 0x02, 0x2B, 0x2D, 0x1F, 0x05, 0x05, 0x04, 0x57, 0x1A,
	0x13, 0x1D, 0x36, 0x5C, 0x3F, 0x74, 0x03, 0x2D, 0x0F, 0x59, 0x28, 0x5B,
	0x03, 0x3A, 0x28, 0x0E, 0x07, 0x19, 0x39, 0x00, 0x08, 0x18, 0x2B, 0x29,
	0x22, 0x1A, 0x1A, 0x2C, 0x17, 0x28, 0x2D, 0x22, 0x50, 0x16, 0x3B, 0x37,
	0x1D, 0x13, 0x3F, 0x58, 0x0D, 0x01, 0x2E, 0x0B, 0x5A, 0x1B, 0x0E, 0x32,
	0x56, 0x27, 0x75, 0x05, 0x28, 0x45, 0x0E, 0x09, 0x0B, 0x33, 0x3A, 0x38,
	0x35, 0x1F, 0x0C, 0x23, 0x3E, 0x3A, 0x0F, 0x0C, 0x07, 0x08, 0x17, 0x3F,
	0x2F, 0x2B, 0x3D, 0x26, 0x01, 0x2B, 0x2B, 0x1E, 0x07, 0x0D, 0x07, 0x2B,
	0x26, 0x2D, 0x0E, 0x2F, 0x3B, 0x20, 0x69, 0x1D, 0x59, 0x1E, 0x2F, 0x17,
	0x07, 0x2E, 0x28, 0x28, 0x2B, 0x38, 0x06, 0x29, 0x1D, 0x3A, 0x1A, 0x14,
	0x00, 0x1C, 0x33, 0x09, 0x11, 0x5C, 0x1F, 0x6D, 0x00, 0x0F, 0x1F, 0x22,
	0x0D, 0x2F, 0x51, 0x34, 0x59, 0x30, 0x0D, 0x51, 0x1F, 0x06, 0x27, 0x1F,
	0x37, 0x09, 0x52, 0x08, 0x3F, 0x0E, 0x0D, 0x2C, 0x07, 0x25, 0x03, 0x08,
	0x21, 0x72, 0x36, 0x0F, 0x5F, 0x25, 0x2F, 0x1E, 0x06, 0x17, 0x29, 0x72,
	0x38, 0x13, 0x5B, 0x3B, 0x14, 0x43, 0x58, 0x28, 0x0F, 0x27, 0x5A, 0x56,
	0x5F, 0x2A, 0x2A, 0x08, 0x37, 0x03, 0x0E, 0x6D, 0x00, 0x30, 0x5D, 0x5A,
	0x33, 0x2E, 0x55, 0x0B, 0x07, 0x11, 0x05, 0x27, 0x3B, 0x3E, 0x25, 0x25,
	0x29, 0x3C, 0x3C, 0x21, 0x29, 0x35, 0x5E, 0x22, 0x33, 0x47, 0x0D, 0x1F,
	0x12, 0x09, 0x1F, 0x16, 0x24, 0x2D, 0x14, 0x3E, 0x13, 0x58, 0x02, 0x2E,
	0x3E, 0x0B, 0x09, 0x5B, 0x01, 0x5B, 0x0E, 0x41, 0x22, 0x0A, 0x21, 0x0A,
	0x2B, 0x19, 0x2F, 0x20, 0x51, 0x06, 0x06, 0x0E, 0x3E, 0x30, 0x00, 0x26,
	0x09, 0x3D, 0x2F, 0x5F, 0x2A, 0x16, 0x58, 0x10, 0x24, 0x00, 0x72, 0x1D,
	0x32, 0x05, 0x12, 0x0C, 0x2A, 0x12, 0x38, 0x07, 0x32, 0x21, 0x30, 0x09,
	0x2F, 0x70, 0x2E, 0x08, 0x01, 0x5C, 0x09, 0x3F, 0x24, 0x1B, 0x26, 0x16,
	0x1C, 0x29, 0x09, 0x1B, 0x05, 0x26, 0x24, 0x01, 0x2E, 0x11, 0x55, 0x37,
	0x05, 0x21, 0x0B, 0x23, 0x51, 0x0A, 0x27, 0x04, 0x5C, 0x0A, 0x26, 0x21,
	0x07, 0x1A, 0x24, 0x19, 0x24, 0x0B, 0x21, 0x23, 0x22, 0x13, 0x04, 0x2E,
	0x52, 0x22, 0x39, 0x76, 0x27, 0x24, 0x38, 0x5F, 0x73, 0x08, 0x54, 0x3F,
	0x06, 0x12, 0x39, 0x16, 0x0B, 0x5E, 0x2C, 0x5C, 0x03, 0x02, 0x44, 0x18,
	0x34, 0x0A, 0x16, 0x1A, 0x21, 0x06, 0x2B, 0x0A, 0x07, 0x6D, 0x5D, 0x0A,
	0x45, 0x59, 0x0E, 0x36, 0x53, 0x2F, 0x21, 0x38, 0x39, 0x05, 0x02, 0x40,
	0x2C, 0x23, 0x19, 0x01, 0x1B, 0x05, 0x1B, 0x17, 0x23, 0x12, 0x1B, 0x59,
	0x2F, 0x07, 0x00, 0x04, 0x3E, 0x35, 0x28, 0x5C, 0x21, 0x19, 0x34, 0x2B,
	0x59, 0x03, 0x0F, 0x03, 0x23, 0x1E, 0x01, 0x21, 0x18, 0x22, 0x1C, 0x73,
	0x28, 0x4A, 0x0D, 0x2A, 0x38, 0x29, 0x0D, 0x04, 0x2E, 0x73, 0x22, 0x0D,
	0x39, 0x0A, 0x11, 0x25, 0x09, 0x1D, 0x09, 0x10, 0x3F, 0x51, 0x3E, 0x2E,
	0x2D, 0x0A, 0x35, 0x1F, 0x39, 0x38, 0x27, 0x3B, 0x3F, 0x12, 0x2B, 0x1E,
	0x53, 0x1C, 0x2D, 0x72, 0x59, 0x15, 0x2F, 0x0D, 0x21, 0x2D, 0x32, 0x41,
	0x1E, 0x06, 0x5C, 0x59, 0x20, 0x3A, 0x1A, 0x1F, 0x0C, 0x37, 0x11, 0x71,
	0x04, 0x10, 0x0A, 0x2E, 0x76, 0x34, 0x31, 0x28, 0x3C, 0x2B, 0x3F, 0x2A,
	0x28, 0x18, 0x27, 0x28, 0x24, 0x1A, 0x5B, 0x21, 0x1F, 0x23, 0x0D, 0x59,
	0x0B, 0x5D, 0x26, 0x23, 0x2C, 0x03, 0x35, 0x58, 0x06, 0x3B, 0x76, 0x2B,
	0x2A, 0x3F, 0x2C, 0x09, 0x0B, 0x2F, 0x2F, 0x29, 0x0E, 0x22, 0x26, 0x22,
	0x08, 0x33, 0x3F, 0x0B, 0x19, 0x12, 0x06, 0x38, 0x11, 0x16, 0x31, 0x72,
	0x28, 0x2A, 0x3A, 0x3E, 0x2E, 0x20, 0x0B, 0x2B, 0x40, 0x0B, 0x1B, 0x51,
	0x1D, 0x38, 0x25, 0x00, 0x22, 0x1E, 0x1B, 0x2A, 0x26, 0x14, 0x21, 0x1F,
	0x76, 0x47, 0x16, 0x04, 0x06, 0x14, 0x2F, 0x2F, 0x2A, 0x23, 0x7A, 0x3E,
	0x04, 0x25, 0x02, 0x1A, 0x27, 0x2A, 0x02, 0x04, 0x11, 0x2D, 0x00, 0x23,
	0x23, 0x11, 0x26, 0x3B, 0x3E, 0x1B, 0x24, 0x07, 0x2D, 0x22, 0x58, 0x75,
	0x28, 0x0E, 0x2B, 0x0D, 0x1B, 0x5A, 0x17, 0x1D, 0x40, 0x13, 0x06, 0x56,
	0x0F, 0x3C, 0x29, 0x1C, 0x10, 0x08, 0x01, 0x30, 0x15, 0x23, 0x2C, 0x29,
	0x0A, 0x28, 0x2F, 0x3B, 0x01, 0x06, 0x3D, 0x3B, 0x3D, 0x32, 0x09, 0x0D,
	0x24, 0x25, 0x20, 0x76, 0x3B, 0x2D, 0x17, 0x04, 0x00, 0x5E, 0x0E, 0x3E,
	0x2E, 0x30, 0x3D, 0x2A, 0x3B, 0x24, 0x35, 0x2A, 0x34, 0x04, 0x19, 0x72,
	0x47, 0x02, 0x3A, 0x24, 0x06, 0x05, 0x08, 0x28, 0x2E, 0x0F, 0x3B, 0x2D,
	0x1E, 0x0A, 0x0E, 0x39, 0x58, 0x22, 0x0C, 0x07, 0x36, 0x15, 0x17, 0x09,
	0x13, 0x06, 0x2E, 0x3D, 0x13, 0x04, 0x05, 0x51, 0x2B, 0x20, 0x10, 0x07,
	0x56, 0x2C, 0x09, 0x13, 0x15, 0x18, 0x0A, 0x2E, 0x2B, 0x35, 0x11, 0x2C,
	0x38, 0x2E, 0x58, 0x38, 0x0D, 0x0F, 0x15, 0x59, 0x20, 0x04, 0x40, 0x06,
	0x15, 0x15, 0x0F, 0x0C, 0x01, 0x54, 0x34, 0x5B, 0x1D, 0x29, 0x36, 0x53,
	0x26, 0x2F, 0x32, 0x0E, 0x2C, 0x1C, 0x22, 0x2E, 0x3E, 0x07, 0x09, 0x3D,
	0x6D, 0x3F, 0x30, 0x03, 0x08, 0x1A, 0x3F, 0x25, 0x28, 0x28, 0x17, 0x3C,
	0x3B, 0x00, 0x31, 0x05, 0x0D, 0x55, 0x1E, 0x04, 0x27, 0x5F, 0x15, 0x1F,
	0x02, 0x34, 0x28, 0x2B, 0x23, 0x3C, 0x17, 0x03, 0x59, 0x1A, 0x26, 0x17,
	0x5C, 0x39, 0x5E, 0x13, 0x11, 0x04, 0x2C, 0x5D, 0x29, 0x04, 0x2B, 0x34,
	0x3C, 0x28, 0x09, 0x3F, 0x3B, 0x1D, 0x2D, 0x0B, 0x00, 0x32, 0x3A, 0x09,
	0x18, 0x5B, 0x56, 0x3E, 0x27, 0x18, 0x26, 0x24, 0x5A, 0x3A, 0x14, 0x2D,
	0x28, 0x3E, 0x59, 0x33, 0x00, 0x11, 0x5A, 0x02, 0x72, 0x5C, 0x06, 0x3C,
	0x31, 0x76, 0x1E, 0x0E, 0x1E, 0x01, 0x1B, 0x24, 0x58, 0x1F, 0x3D, 0x10,
	0x39, 0x12, 0x04, 0x07, 0x2F, 0x1D, 0x00, 0x27, 0x12, 0x27, 0x54, 0x04,
	0x3D, 0x26, 0x0C, 0x2E, 0x22, 0x58, 0x2C, 0x24, 0x01, 0x10, 0x27, 0x26,
	0x37, 0x39, 0x37, 0x27, 0x28, 0x77, 0x1C, 0x18, 0x04, 0x20, 0x35, 0x5F,
	0x00, 0x5A, 0x2A, 0x21, 0x07, 0x19, 0x2D, 0x09, 0x2F, 0x25, 0x03, 0x58,
	0x0C, 0x07, 0x3D, 0x17, 0x01, 0x22, 0x0E, 0x5A, 0x38, 0x3D, 0x07, 0x0C,
	0x38, 0x2C, 0x1D, 0x02, 0x29, 0x21, 0x27, 0x02, 0x26, 0x18, 0x02, 0x30,
	0x2B, 0x1A, 0x08, 0x07, 0x2C, 0x04, 0x32, 0x20, 0x1C, 0x38, 0x2D, 0x08,
	0x10, 0x03, 0x58, 0x56, 0x5B, 0x05, 0x26, 0x11, 0x39, 0x0F, 0x23, 0x01,
	0x3B, 0x03, 0x2E, 0x18, 0x23, 0x08, 0x00, 0x26, 0x3A, 0x39, 0x27, 0x07,
	0x2F, 0x07, 0x26, 0x35, 0x1D, 0x2E, 0x3B, 0x3C, 0x2F, 0x36, 0x28, 0x0C,
	0x03, 0x09, 0x3B, 0x3D, 0x2C, 0x36, 0x0E, 0x03, 0x39, 0x16, 0x19, 0x50,
	0x01, 0x1A, 0x11, 0x1C, 0x08, 0x3A, 0x2F, 0x28, 0x1B, 0x2B, 0x09, 0x2E,
	0x21, 0x5D, 0x00, 0x1A, 0x06, 0x01, 0x06, 0x3B, 0x29, 0x25, 0x08, 0x0F,
	0x36, 0x57, 0x32, 0x70, 0x5E, 0x0C, 0x04, 0x23, 0x0F, 0x0D, 0x53, 0x20,
	0x19, 0x3A, 0x5C, 0x0F, 0x3A, 0x04, 0x14, 0x3B, 0x52, 0x09, 0x2D, 0x13,
	0x22, 0x14, 0x24, 0x5A, 0x73, 0x03, 0x57, 0x22, 0x38, 0x7A, 0x1C, 0x28,
	0x3A, 0x5B, 0x06, 0x25, 0x37, 0x5F, 0x1F, 0x2F, 0x08, 0x3B, 0x2C, 0x59,
	0x0A, 0x23, 0x52, 0x24, 0x58, 0x2A, 0x0B, 0x09, 0x3A, 0x19, 0x01, 0x5E,
	0x17, 0x2F, 0x12, 0x2A, 0x5E, 0x0F, 0x3D, 0x3F, 0x13, 0x23, 0x29, 0x0F,
	0x08, 0x14, 0x26, 0x19, 0x3B, 0x03, 0x09, 0x27, 0x51, 0x27, 0x5E, 0x28,
	0x0E, 0x2E, 0x17, 0x01, 0x28, 0x0F, 0x12, 0x29, 0x0D, 0x14, 0x04, 0x03,
	0x36, 0x1A, 0x77, 0x39, 0x56, 0x0D, 0x3F, 0x72, 0x1C, 0x2F, 0x3C, 0x26,
	0x21, 0x24, 0x20, 0x0F, 0x38, 0x0D, 0x01, 0x32, 0x1F, 0x29, 0x25, 0x14,
	0x32, 0x09, 0x08, 0x32, 0x3D, 0x18, 0x27, 0x29, 0x0E, 0x00, 0x59, 0x59,
	0x06, 0x20, 0x2A, 0x19, 0x05, 0x58, 0x23, 0x15, 0x2E, 0x2A, 0x00, 0x2F,
	0x3B, 0x30, 0x24, 0x52, 0x2A, 0x1C, 0x38, 0x05, 0x26, 0x08, 0x36, 0x15,
	0x16, 0x39, 0x0E, 0x18, 0x0A, 0x1B, 0x5A, 0x1B, 0x03, 0x17, 0x5F, 0x40,
	0x16, 0x02, 0x15, 0x27, 0x24, 0x2B, 0x5B, 0x15, 0x28, 0x3C, 0x72, 0x1B,
	0x0B, 0x01, 0x5E, 0x74, 0x34, 0x37, 0x18, 0x1E, 0x36, 0x1B, 0x10, 0x3F,
	0x26, 0x2F, 0x29, 0x4A, 0x2C, 0x1D, 0x0C, 0x3C, 0x03, 0x38, 0x28, 0x0D,
	0x16, 0x0E, 0x2F, 0x38, 0x34, 0x18, 0x39, 0x29, 0x20, 0x71, 0x3E, 0x24,
	0x09, 0x3F, 0x7A, 0x03, 0x0F, 0x36, 0x39, 0x32, 0x2B, 0x0D, 0x20, 0x0A,
	0x06, 0x3F, 0x19, 0x2A, 0x40, 0x72, 0x36, 0x28, 0x29, 0x5B, 0x31, 0x1C,
	0x2E, 0x21, 0x26, 0x27, 0x23, 0x11, 0x05, 0x13, 0x74, 0x38, 0x30, 0x00,
	0x21, 0x32, 0x02, 0x54, 0x03, 0x5A, 0x34, 0x1D, 0x2C, 0x2A, 0x0C, 0x73,
	0x2B, 0x0C, 0x01, 0x0C, 0x14, 0x58, 0x59, 0x19, 0x3D, 0x76, 0x2A, 0x17,
	0x3C, 0x58, 0x34, 0x0E, 0x36, 0x2D, 0x0C, 0x37, 0x0E, 0x20, 0x5C, 0x2A,
	0x69, 0x14, 0x52, 0x45, 0x11, 0x76, 0x23, 0x07, 0x34, 0x58, 0x01, 0x0B,
	0x11, 0x5D, 0x40, 0x14, 0x34, 0x57, 0x5C, 0x2A, 0x69, 0x14, 0x52, 0x45,
	0x31, 0x35, 0x38, 0x59, 0x27, 0x07, 0x14, 0x5C, 0x37, 0x22, 0x1B, 0x1B,
	0x34, 0x0B, 0x08, 0x0F, 0x25, 0x2D, 0x12, 0x38, 0x0E, 0x25, 0x36, 0x39,
	0x5F, 0x0F, 0x20, 0x1A, 0x56, 0x0C, 0x40, 0x3A, 0x20, 0x35, 0x25, 0x18,
	0x69, 0x0A, 0x17, 0x1C, 0x01, 0x15, 0x1A, 0x09, 0x5B, 0x0E, 0x31, 0x1C,
	0x22, 0x34, 0x3F, 0x15, 0x0F, 0x4E, 0x07, 0x52, 0x6D, 0x08, 0x54, 0x45,
	0x09, 0x6D, 0x47, 0x2D, 0x20, 0x03, 0x27, 0x3F, 0x4E, 0x04, 0x5C, 0x75,
	0x1F, 0x30, 0x22, 0x5F, 0x0B, 0x15, 0x25, 0x1E, 0x0F, 0x26, 0x59, 0x02,
	0x56, 0x02, 0x0E, 0x16, 0x12, 0x18, 0x26, 0x13, 0x0A, 0x09, 0x2B, 0x20,
	0x7A, 0x3D, 0x24, 0x1F, 0x28, 0x2E, 0x1B, 0x2A, 0x2C, 0x32, 0x15, 0x3E,
	0x09, 0x3F, 0x06, 0x04, 0x07, 0x12, 0x24, 0x03, 0x2A, 0x38, 0x0C, 0x28,
	0x28, 0x35, 0x03, 0x2D, 0x2D, 0x5B, 0x31, 0x27, 0x05, 0x16, 0x38, 0x15,
	0x2A, 0x09, 0x5A, 0x19, 0x0E, 0x2F, 0x12, 0x1D, 0x27, 0x74, 0x1B, 0x0E,
	0x08, 0x2D, 0x3A, 0x35, 0x36, 0x3F, 0x02, 0x09, 0x5E, 0x32, 0x3C, 0x12,
	0x03, 0x08, 0x08, 0x16, 0x1D, 0x05, 0x14, 0x54, 0x16, 0x33, 0x08, 0x39,
	0x13, 0x28, 0x3D, 0x31, 0x3B, 0x26, 0x16, 0x38, 0x38, 0x2F, 0x14, 0x5C,
	0x20, 0x37, 0x35, 0x39, 0x21, 0x13, 0x15, 0x5B, 0x27, 0x3E, 0x18, 0x17,
	0x2F, 0x55, 0x01, 0x01, 0x2B, 0x05, 0x2E, 0x22, 0x2E, 0x76, 0x03, 0x0D,
	0x16, 0x08, 0x0D, 0x27, 0x12, 0x5A, 0x18, 0x2C, 0x2A, 0x04, 0x0D, 0x3D,
	0x04, 0x14, 0x00, 0x36, 0x2D, 0x0D, 0x54, 0x0E, 0x22, 0x02, 0x72, 0x47,
	0x37, 0x02, 0x13, 0x15, 0x06, 0x24, 0x1E, 0x21, 0x36, 0x2D, 0x56, 0x07,
	0x07, 0x74, 0x58, 0x55, 0x1A, 0x1A, 0x08, 0x1F, 0x33, 0x08, 0x06, 0x09,
	0x14, 0x18, 0x1D, 0x1A, 0x14, 0x5A, 0x2F, 0x56, 0x1C, 0x71, 0x14, 0x04,
	0x3E, 0x01, 0x6D, 0x0A, 0x2B, 0x38, 0x40, 0x13, 0x24, 0x54, 0x05, 0x1D,
	0x3B, 0x0F, 0x4E, 0x21, 0x11, 0x7A, 0x02, 0x31, 0x17, 0x12, 0x6D, 0x26,
	0x2D, 0x56, 0x5B, 0x34, 0x15, 0x57, 0x41, 0x22, 0x30, 0x54, 0x19, 0x26,
	0x29, 0x1B, 0x35, 0x27, 0x18, 0x2A, 0x08, 0x47, 0x06, 0x3B, 0x1E, 0x00,
	0x03, 0x22, 0x2D, 0x12, 0x13, 0x2A, 0x2A, 0x3F, 0x33, 0x18, 0x2E, 0x35,
	0x05, 0x2D, 0x26, 0x3D, 0x34, 0x02, 0x29, 0x23, 0x39, 0x27, 0x34, 0x3A,
	0x17, 0x3A, 0x23, 0x34, 0x0C, 0x03, 0x03, 0x2F, 0x2D, 0x58, 0x2F, 0x2A,
	0x4E, 0x2B, 0x21, 0x18, 0x2F, 0x32, 0x3D, 0x2D, 0x70, 0x3B, 0x23, 0x41,
	0x23, 0x2E, 0x04, 0x07, 0x2D, 0x1B, 0x18, 0x34, 0x38, 0x25, 0x1D, 0x1A,
	0x2B, 0x2A, 0x59, 0x03, 0x30, 0x09, 0x26, 0x18, 0x08, 0x14, 0x07, 0x0B,
	0x39, 0x29, 0x0D, 0x59, 0x33, 0x1C, 0x22, 0x2F, 0x09, 0x51, 0x5D, 0x24,
	0x2F, 0x1E, 0x16, 0x5F, 0x21, 0x15, 0x18, 0x2A, 0x5F, 0x5E, 0x11, 0x18,
	0x10, 0x38, 0x03, 0x16, 0x19, 0x30, 0x37, 0x3D, 0x05, 0x3E, 0x03, 0x16,
	0x02, 0x34, 0x04, 0x27, 0x22, 0x00, 0x15, 0x2F, 0x0E, 0x1D, 0x0C, 0x2B,
	0x3F, 0x37, 0x28, 0x59, 0x17, 0x39, 0x54, 0x3C, 0x33, 0x2E, 0x2A, 0x2B,
	0x2B, 0x0E, 0x08, 0x1E, 0x51, 0x22, 0x5C, 0x11, 0x15, 0x14, 0x3E, 0x07,
	0x0D, 0x09, 0x36, 0x5B, 0x5E, 0x12, 0x5D, 0x52, 0x25, 0x1E, 0x6D, 0x43,
	0x07, 0x22, 0x25, 0x05, 0x1F, 0x0B, 0x36, 0x5A, 0x04, 0x2F, 0x17, 0x58,
	0x0F, 0x18, 0x23, 0x2F, 0x5B, 0x44, 0x23, 0x5D, 0x57, 0x2A, 0x0E, 0x28,
	0x55, 0x00, 0x5C, 0x1A, 0x7B, 0x24, 0x58, 0x18, 0x44, 0x74, 0x19, 0x52,
	0x5F, 0x0C, 0x2B, 0x1A, 0x11, 0x3B, 0x01, 0x13, 0x00, 0x32, 0x05, 0x5C,
	0x28, 0x5B, 0x2C, 0x0C, 0x0C, 0x03, 0x3B, 0x24, 0x3A, 0x23, 0x35, 0x07,
	0x14, 0x5A, 0x06, 0x00, 0x38, 0x20, 0x45, 0x1D, 0x01, 0x5A, 0x1B, 0x1E,
	0x23, 0x10, 0x06, 0x2A, 0x0D, 0x40, 0x6D, 0x0B, 0x18, 0x22, 0x11, 0x31,
	0x16, 0x13, 0x20, 0x21, 0x2E, 0x01, 0x00, 0x05, 0x02, 0x0E, 0x1A, 0x29,
	0x5A, 0x5A, 0x34, 0x22, 0x08, 0x3A, 0x2C, 0x35, 0x2B, 0x54, 0x3B, 0x3C,
	0x29, 0x55, 0x23, 0x57, 0x06, 0x04, 0x22, 0x0F, 0x03, 0x53, 0x76, 0x23,
	0x31, 0x24, 0x1F, 0x76, 0x47, 0x07, 0x56, 0x0C, 0x69, 0x5A, 0x0E, 0x3F,
	0x21, 0x6D, 0x2E, 0x50, 0x06, 0x5C, 0x6D, 0x58, 0x2F, 0x36, 0x1A, 0x7A,
	0x55, 0x2B, 0x5F, 0x25, 0x17, 0x01, 0x2B, 0x5E, 0x0D, 0x03, 0x14, 0x24,
	0x04, 0x3E, 0x36, 0x26, 0x15, 0x0F, 0x2D, 0x1A, 0x1F, 0x03, 0x3D, 0x39,
	0x3B, 0x23, 0x54, 0x28, 0x1C, 0x1A, 0x3A, 0x37, 0x56, 0x40, 0x0D, 0x21,
	0x27, 0x08, 0x5B, 0x10, 0x1A, 0x12, 0x21, 0x0C, 0x07, 0x35, 0x31, 0x18,
	0x2C, 0x18, 0x26, 0x00, 0x03, 0x00, 0x2F, 0x1C, 0x2A, 0x08, 0x2E, 0x7A,
	0x47, 0x0A, 0x57, 0x2C, 0x01, 0x1E, 0x55, 0x0D, 0x2E, 0x7A, 0x0A, 0x18,
	0x2B, 0x1E, 0x07, 0x15, 0x0F, 0x57, 0x39, 0x11, 0x1E, 0x1B, 0x1E, 0x28,
	0x07, 0x5A, 0x33, 0x03, 0x0E, 0x25, 0x26, 0x02, 0x5D, 0x38, 0x2F, 0x1C,
	0x10, 0x0F, 0x00, 0x38, 0x39, 0x2A, 0x39, 0x04, 0x32, 0x1F, 0x0D, 0x38,
	0x26, 0x14, 0x3F, 0x0B, 0x04, 0x53, 0x2C, 0x3B, 0x28, 0x27, 0x3C, 0x31,
	0x18, 0x33, 0x3D, 0x23, 0x05, 0x3E, 0x17, 0x3B, 0x5E, 0x0B, 0x0A, 0x34,
	0x5F, 0x24, 0x0E, 0x1B, 0x0C, 0x1F, 0x21, 0x0B, 0x3F, 0x59, 0x1D, 0x2C,
	0x2C, 0x27, 0x02, 0x20, 0x20, 0x26, 0x3A, 0x06, 0x29, 0x20, 0x29, 0x19,
	0x12, 0x19, 0x3B, 0x34, 0x39, 0x28, 0x02, 0x5F, 0x18, 0x3D, 0x29, 0x1D,
	0x25, 0x3A, 0x2A, 0x02, 0x39, 0x12, 0x20, 0x2F, 0x3B, 0x3A, 0x5D, 0x74,
	0x06, 0x4E, 0x2F, 0x19, 0x34, 0x03, 0x31, 0x16, 0x00, 0x75, 0x54, 0x33,
	0x0D, 0x28, 0x35, 0x07, 0x2F, 0x20, 0x29, 0x16, 0x26, 0x29, 0x3A, 0x58,
	0x7A, 0x0A, 0x30, 0x27, 0x52, 0x24, 0x08, 0x0A, 0x0D, 0x1C, 0x0E, 0x34,
	0x55, 0x2C, 0x29, 0x24, 0x3A, 0x52, 0x57, 0x39, 0x31, 0x27, 0x04, 0x5D,
	0x12, 0x0F, 0x22, 0x35, 0x5A, 0x29, 0x2C, 0x03, 0x55, 0x3C, 0x05, 0x2D,
	0x5F, 0x06, 0x0D, 0x39, 0x30, 0x2A, 0x0B, 0x2D, 0x3C, 0x30, 0x34, 0x28,
	0x5C, 0x19, 0x15, 0x54, 0x23, 0x2D, 0x27, 0x71, 0x03, 0x2C, 0x2F, 0x1C,
	0x38, 0x47, 0x20, 0x3F, 0x22, 0x16, 0x1F, 0x26, 0x38, 0x33, 0x37, 0x21,
	0x0C, 0x1A, 0x3F, 0x14, 0x1D, 0x15, 0x3F, 0x52, 0x12, 0x25, 0x34, 0x06,
	0x22, 0x2B, 0x55, 0x39, 0x08, 0x12, 0x07, 0x3B, 0x23, 0x3D, 0x20, 0x34,
	0x03, 0x26, 0x2D, 0x39, 0x36, 0x5B, 0x59, 0x59, 0x3E, 0x37, 0x0F, 0x0C,
	0x25, 0x29, 0x16, 0x58, 0x4A, 0x5A, 0x09, 0x25, 0x59, 0x28, 0x3C, 0x22,
	0x2D, 0x5F, 0x0E, 0x06, 0x1D, 0x24, 0x14, 0x05, 0x18, 0x0E, 0x2F, 0x54,
	0x09, 0x2D, 0x2C, 0x37, 0x43, 0x17, 0x5B, 0x22, 0x31, 0x5C, 0x0E, 0x04,
	0x22, 0x01, 0x0B, 0x12, 0x2F, 0x06, 0x2F, 0x14, 0x58, 0x04, 0x5B, 0x06,
	0x0B, 0x0E, 0x22, 0x5C, 0x2B, 0x2D, 0x2B, 0x56, 0x03, 0x13, 0x2B, 0x14,
	0x27, 0x0E, 0x76, 0x47, 0x35, 0x2F, 0x3F, 0x36, 0x27, 0x06, 0x3B, 0x1D,
	0x37, 0x21, 0x55, 0x3F, 0x1E, 0x13, 0x0F, 0x28, 0x3C, 0x20, 0x74, 0x2E,
	0x29, 0x07, 0x20, 0x71, 0x35, 0x2F, 0x0A, 0x2A, 0x17, 0x23, 0x11, 0x01,
	0x01, 0x71, 0x38, 0x10, 0x5F, 0x1E, 0x28, 0x1F, 0x06, 0x26, 0x3F, 0x30,
	0x5D, 0x09, 0x2F, 0x2C, 0x1B, 0x3F, 0x2E, 0x28, 0x38, 0x07, 0x55, 0x2B,
	0x14, 0x0F, 0x17, 0x43, 0x0D, 0x25, 0x3C, 0x05, 0x5A, 0x0D, 0x3B, 0x0F,
	0x26, 0x02, 0x37, 0x5D, 0x2F, 0x35, 0x5C, 0x28, 0x57, 0x33, 0x21, 0x22,
	0x59, 0x3C, 0x3A, 0x04, 0x04, 0x38, 0x34, 0x5F, 0x00, 0x43, 0x0A, 0x29,
	0x0E, 0x2D, 0x18, 0x02, 0x09, 0x12, 0x07, 0x26, 0x07, 0x34, 0x32, 0x06,
	0x0B, 0x0E, 0x3E, 0x53, 0x25, 0x5B, 0x19, 0x2A, 0x3B, 0x17, 0x3B, 0x09,
	0x3F, 0x05, 0x35, 0x35, 0x32, 0x1B, 0x1E, 0x08, 0x28, 0x2A, 0x01, 0x24,
	0x27, 0x1B, 0x11, 0x56, 0x1A, 0x3A, 0x5C, 0x53, 0x1C, 0x2F, 0x33, 0x21,
	0x59, 0x41, 0x0D, 0x71, 0x08, 0x20, 0x36, 0x38, 0x2B, 0x26, 0x37, 0x05,
	0x1A, 0x0C, 0x2F, 0x29, 0x0D, 0x39, 0x0D, 0x1D, 0x1B, 0x58, 0x04, 0x07,
	0x3F, 0x2C, 0x2C, 0x0D, 0x26, 0x04, 0x30, 0x34, 0x18, 0x70, 0x03, 0x17,
	0x25, 0x25, 0x10, 0x22, 0x35, 0x04, 0x0E, 0x2D, 0x1E, 0x09, 0x5E, 0x00,
	0x13, 0x2D, 0x53, 0x1C, 0x20, 0x35, 0x3C, 0x03, 0x07, 0x2D, 0x70, 0x26,
	0x29, 0x07, 0x20, 0x2A, 0x38, 0x50, 0x2F, 0x1C, 0x36, 0x25, 0x2D, 0x3F,
	0x3A, 0x12, 0x0F, 0x30, 0x5D, 0x5D, 0x00, 0x2D, 0x50, 0x24, 0x03, 0x75,
	0x22, 0x2F, 0x09, 0x11, 0x08, 0x28, 0x30, 0x5A, 0x3E, 0x0B, 0x04, 0x2C,
	0x39, 0x27, 0x76, 0x20, 0x22, 0x09, 0x5B, 0x15, 0x55, 0x30, 0x01, 0x2D,
	0x0A, 0x43, 0x17, 0x59, 0x29, 0x34, 0x05, 0x26, 0x01, 0x28, 0x23, 0x1F,
	0x17, 0x27, 0x24, 0x7A, 0x3D, 0x12, 0x24, 0x0F, 0x25, 0x5B, 0x27, 0x14,
	0x3B, 0x0E, 0x5C, 0x59, 0x01, 0x31, 0x08, 0x14, 0x51, 0x0A, 0x5B, 0x7A,
	0x2D, 0x1B, 0x5C, 0x52, 0x24, 0x22, 0x53, 0x06, 0x18, 0x23, 0x2F, 0x0C,
	0x38, 0x0A, 0x30, 0x47, 0x56, 0x09, 0x20, 0x2F, 0x2E, 0x3B, 0x06, 0x3C,
	0x29, 0x0F, 0x26, 0x0B, 0x00, 0x05, 0x3A, 0x20, 0x05, 0x22, 0x27, 0x1A,
	0x37, 0x16, 0x44, 0x2D, 0x0D, 0x33, 0x16, 0x05, 0x69, 0x3D, 0x00, 0x58,
	0x0E, 0x71, 0x05, 0x57, 0x01, 0x40, 0x18, 0x3A, 0x13, 0x29, 0x52, 0x25,
	0x05, 0x2A, 0x0B, 0x58, 0x18, 0x5B, 0x25, 0x27, 0x1C, 0x35, 0x18, 0x08,
	0x5E, 0x26, 0x71, 0x22, 0x34, 0x5A, 0x03, 0x23, 0x3A, 0x23, 0x5E, 0x3B,
	0x07, 0x03, 0x32, 0x27, 0x33, 0x0E, 0x5D, 0x25, 0x3B, 0x3E, 0x36, 0x3B,
	0x17, 0x37, 0x32, 0x04, 0x47, 0x39, 0x1E, 0x0C, 0x34, 0x55, 0x2F, 0x1A,
	0x58, 0x26, 0x34, 0x25, 0x27, 0x13, 0x28, 0x14, 0x36, 0x20, 0x09, 0x75,
	0x2E, 0x55, 0x39, 0x27, 0x24, 0x27, 0x29, 0x0B, 0x5F, 0x17, 0x55, 0x20,
	0x3C, 0x58, 0x36, 0x0F, 0x24, 0x56, 0x02, 0x31, 0x00, 0x12, 0x20, 0x24,
	0x3B, 0x2A, 0x16, 0x5B, 0x3C, 0x14, 0x2F, 0x29, 0x3E, 0x20, 0x07, 0x55,
	0x55, 0x0C, 0x3F, 0x26, 0x5A, 0x30, 0x1E, 0x1D, 0x14, 0x0D, 0x50, 0x0F,
	0x03, 0x01, 0x24, 0x23, 0x27, 0x2E, 0x03, 0x18, 0x15, 0x29, 0x0A, 0x71,
	0x26, 0x29, 0x2C, 0x3C, 0x31, 0x21, 0x06, 0x18, 0x26, 0x01, 0x0B, 0x59,
	0x2B, 0x2D, 0x35, 0x0B, 0x16, 0x2B, 0x3E, 0x10, 0x19, 0x0E, 0x28, 0x1A,
	0x29, 0x22, 0x20, 0x20, 0x3C, 0x20, 0x2D, 0x57, 0x05, 0x20, 0x6D, 0x3D,
	0x50, 0x0A, 0x44, 0x1A, 0x23, 0x58, 0x2A, 0x3F, 0x25, 0x15, 0x55, 0x1D,
	0x00, 0x3A, 0x36, 0x14, 0x07, 0x22, 0x30, 0x3B, 0x2B, 0x05, 0x38, 0x15,
	0x34, 0x2D, 0x0D, 0x21, 0x1A, 0x34, 0x53, 0x56, 0x3E, 0x00, 0x1F, 0x14,
	0x5B, 0x40, 0x76, 0x0A, 0x55, 0x01, 0x2C, 0x31, 0x19, 0x2B, 0x16, 0x09,
	0x01, 0x2B, 0x10, 0x1C, 0x33, 0x01, 0x28, 0x14, 0x17, 0x24, 0x03, 0x3B,
	0x55, 0x27, 0x1D, 0x23, 0x1F, 0x37, 0x3F, 0x53, 0x27, 0x03, 0x39, 0x2D,
	0x5D, 0x00, 0x29, 0x00, 0x2D, 0x25, 0x71, 0x2D, 0x29, 0x59, 0x3D, 0x2C,
	0x19, 0x33, 0x5F, 0x33, 0x28, 0x3E, 0x02, 0x57, 0x52, 0x07, 0x2D, 0x37,
	0x2D, 0x3A, 0x0D, 0x3E, 0x05, 0x3A, 0x3D, 0x0A, 0x09, 0x02, 0x28, 0x2A,
	0x77, 0x25, 0x0D, 0x1D, 0x3C, 0x08, 0x5C, 0x0D, 0x3F, 0x04, 0x03, 0x5B,
	0x0E, 0x1F, 0x1E, 0x20, 0x29, 0x2F, 0x02, 0x12, 0x75, 0x0A, 0x2D, 0x16,
	0x1B, 0x11, 0x1A, 0x39, 0x17, 0x13, 0x26, 0x0F, 0x3B, 0x1F, 0x0F, 0x17,
	0x22, 0x2F, 0x37, 0x03, 0x12, 0x1A, 0x04, 0x3F, 0x07, 0x73, 0x09, 0x16,
	0x1E, 0x5D, 0x21, 0x2D, 0x05, 0x39, 0x2F, 0x2C, 0x29, 0x22, 0x24, 0x12,
	0x76, 0x02, 0x05, 0x5E, 0x08, 0x31, 0x3F, 0x26, 0x3F, 0x09, 0x31, 0x20,
	0x25, 0x2C, 0x2E, 0x2B, 0x47, 0x57, 0x1C, 0x2F, 0x71, 0x18, 0x23, 0x29,
	0x0C, 0x70, 0x3B, 0x25, 0x1E, 0x1B, 0x03, 0x36, 0x58, 0x26, 0x12, 0x2A,
	0x3B, 0x23, 0x5C, 0x5E, 0x0B, 0x5E, 0x27, 0x01, 0x04, 0x0C, 0x16, 0x4E,
	0x41, 0x00, 0x0A, 0x3D, 0x34, 0x25, 0x2C, 0x00, 0x47, 0x30, 0x34, 0x2A,
	0x33, 0x5F, 0x00, 0x01, 0x3F, 0x13, 0x18, 0x10, 0x23, 0x25, 0x2A, 0x38,
	0x0E, 0x0A, 0x31, 0x08, 0x09, 0x3B, 0x16, 0x59, 0x7B, 0x54, 0x2C, 0x58,
	0x18, 0x2C, 0x0D, 0x23, 0x3E, 0x0A, 0x1A, 0x3D, 0x56, 0x23, 0x11, 0x14,
	0x28, 0x2E, 0x05, 0x01, 0x7A, 0x3C, 0x35, 0x5D, 0x2D, 0x03, 0x1C, 0x0D,
	0x58, 0x3A, 0x2F, 0x3E, 0x28, 0x41, 0x08, 0x35, 0x18, 0x0E, 0x3B, 0x1D,
	0x21, 0x19, 0x12, 0x04, 0x2E, 0x29, 0x3D, 0x24, 0x2C, 0x38, 0x0F, 0x02,
	0x03, 0x09, 0x08, 0x08, 0x2E, 0x0F, 0x20, 0x0C, 0x7B, 0x27, 0x38, 0x59,
	0x03, 0x3B, 0x0B, 0x0A, 0x3D, 0x29, 0x13, 0x2B, 0x07, 0x0F, 0x03, 0x0E,
	0x24, 0x32, 0x1E, 0x0E, 0x35, 0x39, 0x24, 0x2C, 0x1F, 0x08, 0x26, 0x1B,
	0x04, 0x3E, 0x33, 0x15, 0x24, 0x5A, 0x04, 0x13, 0x2E, 0x06, 0x01, 0x03,
	0x74, 0x1F, 0x0E, 0x17, 0x0C, 0x38, 0x59, 0x27, 0x0D, 0x2F, 0x2D, 0x2D,
	0x57, 0x5C, 0x38, 0x04, 0x19, 0x0F, 0x28, 0x19, 0x00, 0x59, 0x28, 0x3E,
	0x3E, 0x26, 0x20, 0x0E, 0x36, 0x1A, 0x0D, 0x2B, 0x55, 0x00, 0x2A, 0x12,
	0x1C, 0x37, 0x5A, 0x04, 0x07, 0x3C, 0x10, 0x2B, 0x0E, 0x30, 0x01, 0x09,
	0x00, 0x18, 0x2D, 0x18, 0x18, 0x56, 0x2C, 0x36, 0x38, 0x55, 0x07, 0x18,
	0x12, 0x43, 0x0D, 0x29, 0x0C, 0x09, 0x22, 0x02, 0x1B, 0x20, 0x2E, 0x5A,
	0x14, 0x5A, 0x09, 0x76, 0x3D, 0x24, 0x26, 0x18, 0x7A, 0x0D, 0x0D, 0x22,
	0x02, 0x04, 0x14, 0x13, 0x3E, 0x24, 0x25, 0x0B, 0x2E, 0x45, 0x03, 0x15,
	0x5C, 0x51, 0x26, 0x00, 0x30, 0x1C, 0x19, 0x08, 0x29, 0x71, 0x1F, 0x0F,
	0x1C, 0x1C, 0x00, 0x34, 0x0A, 0x0C, 0x1E, 0x12, 0x27, 0x58, 0x3F, 0x0D,
	0x7A, 0x00, 0x20, 0x45, 0x09, 0x0C, 0x47, 0x11, 0x23, 0x40, 0x37, 0x1B,
	0x3B, 0x57, 0x33, 0x2A, 0x21, 0x29, 0x1D, 0x3B, 0x0E, 0x5E, 0x09, 0x1C,
	0x23, 0x33, 0x24, 0x51, 0x03, 0x28, 0x31, 0x0A, 0x20, 0x26, 0x13, 0x25,
	0x3D, 0x23, 0x24, 0x5F, 0x0B, 0x2F, 0x58, 0x5C, 0x26, 0x2A, 0x2B, 0x30,
	0x3C, 0x06, 0x71, 0x18, 0x1B, 0x1C, 0x18, 0x0D, 0x3E, 0x36, 0x59, 0x3F,
	0x7A, 0x5A, 0x0C, 0x03, 0x12, 0x16, 0x1D, 0x11, 0x45, 0x58, 0x0B, 0x23,
	0x30, 0x1E, 0x2E, 0x17, 0x5C, 0x39, 0x1E, 0x3D, 0x2B, 0x15, 0x38, 0x41,
	0x5F, 0x2E, 0x0A, 0x15, 0x2D, 0x2F, 0x72, 0x05, 0x55, 0x3B, 0x09, 0x2D,
	0x5A, 0x4A, 0x05, 0x24, 0x30, 0x1A, 0x04, 0x18, 0x05, 0x2B, 0x22, 0x15,
	0x3B, 0x31, 0x14, 0x2B, 0x20, 0x2B, 0x0E, 0x28, 0x39, 0x16, 0x0A, 0x5C,
	0x77, 0x3F, 0x30, 0x2D, 0x1A, 0x3B, 0x07, 0x0E, 0x24, 0x13, 0x04, 0x39,
	0x56, 0x08, 0x1C, 0x15, 0x5B, 0x09, 0x18, 0x02, 0x25, 0x54, 0x05, 0x5F,
	0x21, 0x05, 0x2E, 0x27, 0x57, 0x0C, 0x7B, 0x5F, 0x56, 0x3F, 0x26, 0x36,
	0x2B, 0x51, 0x59, 0x12, 0x0F, 0x3C, 0x14, 0x2F, 0x06, 0x2A, 0x38, 0x23,
	0x23, 0x22, 0x00, 0x5A, 0x12, 0x5C, 0x1A, 0x1B, 0x24, 0x12, 0x3E, 0x1C,
	0x21, 0x23, 0x13, 0x18, 0x2C, 0x1B, 0x05, 0x22, 0x39, 0x3C, 0x71, 0x22,
	0x19, 0x57, 0x08, 0x30, 0x1C, 0x20, 0x23, 0x38, 0x14, 0x06, 0x27, 0x57,
	0x3B, 0x24, 0x2A, 0x06, 0x29, 0x13, 0x07, 0x2F, 0x0A, 0x17, 0x00, 0x2F,
	0x1E, 0x51, 0x2F, 0x3B, 0x04, 0x21, 0x2A, 0x34, 0x2D, 0x03, 0x3D, 0x24,
	0x06, 0x38, 0x2B, 0x2B, 0x2D, 0x36, 0x12, 0x70, 0x3D, 0x2A, 0x29, 0x18,
	0x17, 0x5A, 0x02, 0x1C, 0x2F, 0x08, 0x01, 0x18, 0x5B, 0x04, 0x2C, 0x2F,
	0x00, 0x04, 0x11, 0x36, 0x05, 0x02, 0x25, 0x2F, 0x24, 0x39, 0x2C, 0x56,
	0x3E, 0x16, 0x04, 0x0F, 0x29, 0x0C, 0x14, 0x43, 0x2E, 0x01, 0x01, 0x01,
	0x0A, 0x27, 0x5F, 0x2D, 0x72, 0x20, 0x59, 0x04, 0x1A, 0x2D, 0x58, 0x24,
	0x2C, 0x1E, 0x0A, 0x14, 0x37, 0x45, 0x2F, 0x33, 0x2B, 0x4A, 0x19, 0x20,
	0x18, 0x39, 0x05, 0x57, 0x0A, 0x32, 0x5A, 0x23, 0x17, 0x00, 0x74, 0x15,
	0x07, 0x0F, 0x1D, 0x20, 0x5E, 0x2B, 0x1B, 0x59, 0x07, 0x0A, 0x36, 0x1C,
	0x12, 0x1A, 0x1C, 0x3B, 0x17, 0x40, 0x2A, 0x0A, 0x05, 0x37, 0x0C, 0x32,
	0x29, 0x29, 0x37, 0x0D, 0x05, 0x1D, 0x25, 0x0D, 0x53, 0x24, 0x5E, 0x25,
	0x03, 0x29, 0x2F, 0x23, 0x24, 0x2F, 0x58, 0x29, 0x08, 0x11, 0x19, 0x22,
	0x26, 0x14, 0x58, 0x18, 0x25, 0x3B, 0x38, 0x08, 0x05, 0x1A, 0x06, 0x26,
	0x33, 0x5B, 0x23, 0x21, 0x0F, 0x12, 0x06, 0x5D, 0x12, 0x2B, 0x50, 0x3F,
	0x07, 0x0A, 0x25, 0x52, 0x37, 0x00, 0x1B, 0x28, 0x2E, 0x3E, 0x58, 0x28,
	0x1B, 0x58, 0x28, 0x3D, 0x2A, 0x59, 0x0F, 0x5B, 0x23, 0x16, 0x06, 0x34,
	0x19, 0x5A, 0x24, 0x3B, 0x0A, 0x5C, 0x2F, 0x01, 0x2D, 0x03, 0x5E, 0x58,
	0x32, 0x07, 0x10, 0x02, 0x25, 0x7A, 0x1A, 0x14, 0x5C, 0x21, 0x32, 0x54,
	0x28, 0x2D, 0x1E, 0x32, 0x01, 0x29, 0x39, 0x06, 0x25, 0x28, 0x0C, 0x20,
	0x20, 0x03, 0x14, 0x39, 0x0A, 0x20, 0x2A, 0x2D, 0x20, 0x24, 0x5B, 0x69,
	0x06, 0x0B, 0x38, 0x05, 0x25, 0x09, 0x11, 0x2A, 0x53, 0x21, 0x15, 0x0D,
	0x2F, 0x09, 0x74, 0x2B, 0x55, 0x02, 0x1C, 0x23, 0x5B, 0x22, 0x2A, 0x0E,
	0x3B, 0x2F, 0x59, 0x20, 0x33, 0x0B, 0x3C, 0x23, 0x22, 0x2F, 0x35, 0x2A,
	0x55, 0x21, 0x5F, 0x0E, 0x1F, 0x25, 0x1B, 0x32, 0x74, 0x1B, 0x20, 0x5C,
	0x5E, 0x27, 0x38, 0x26, 0x3A, 0x3B, 0x36, 0x1C, 0x2C, 0x09, 0x20, 0x71,
	0x34, 0x57, 0x1E, 0x1A, 0x71, 0x5C, 0x51, 0x37, 0x5C, 0x2B, 0x1C, 0x06,
	0x1E, 0x1E, 0x72, 0x5C, 0x30, 0x34, 0x1E, 0x2A, 0x06, 0x10, 0x45, 0x5B,
	0x0D, 0x2E, 0x02, 0x59, 0x03, 0x37, 0x1E, 0x51, 0x0C, 0x44, 0x0E, 0x3D,
	0x06, 0x3B, 0x23, 0x15, 0x00, 0x2C, 0x1B, 0x20, 0x11, 0x14, 0x18, 0x5A,
	0x1D, 0x04, 0x29, 0x35, 0x5E, 0x39, 0x7B, 0x3B, 0x57, 0x20, 0x2A, 0x18,
	0x1E, 0x0E, 0x0B, 0x04, 0x2F, 0x2A, 0x35, 0x56, 0x40, 0x1B, 0x22, 0x09,
	0x18, 0x28, 0x32, 0x23, 0x32, 0x56, 0x23, 0x08, 0x1E, 0x11, 0x38, 0x22,
	0x13, 0x1B, 0x34, 0x06, 0x1D, 0x76, 0x16, 0x08, 0x25, 0x39, 0x28, 0x23,
	0x09, 0x34, 0x0E, 0x2A, 0x3C, 0x26, 0x39, 0x08, 0x0C, 0x5C, 0x59, 0x5B,
	0x0A, 0x11, 0x2E, 0x50, 0x56, 0x2F, 0x0F, 0x29, 0x28, 0x01, 0x00, 0x17,
	0x16, 0x26, 0x16, 0x05, 0x70, 0x2D, 0x00, 0x1B, 0x1C, 0x0C, 0x3F, 0x36,
	0x58, 0x02, 0x0D, 0x5C, 0x32, 0x16, 0x52, 0x6D, 0x5D, 0x16, 0x0C, 0x26,
	0x32, 0x19, 0x17, 0x36, 0x58, 0x3A, 0x0F, 0x57, 0x06, 0x1C, 0x28, 0x36,
	0x03, 0x3F, 0x2A, 0x15, 0x23, 0x20, 0x56, 0x3C, 0x3A, 0x54, 0x02, 0x0D,
	0x23, 0x27, 0x39, 0x2F, 0x2C, 0x27, 0x72, 0x0F, 0x4A, 0x02, 0x1B, 0x1B,
	0x2D, 0x51, 0x0B, 0x0D, 0x2D, 0x5F, 0x51, 0x36, 0x44, 0x2F, 0x1C, 0x35,
	0x0B, 0x08, 0x3B, 0x15, 0x19, 0x06, 0x1B, 0x2C, 0x35, 0x25, 0x0B, 0x33,
	0x0B, 0x34, 0x2E, 0x3B, 0x5A, 0x76, 0x0E, 0x4A, 0x36, 0x5C, 0x25, 0x3E,
	0x33, 0x1D, 0x02, 0x35, 0x1F, 0x33, 0x28, 0x39, 0x71, 0x58, 0x25, 0x3D,
	0x25, 0x7B, 0x3B, 0x52, 0x5E, 0x2F, 0x27, 0x01, 0x17, 0x58, 0x1F, 0x25,
	0x04, 0x32, 0x07, 0x1F, 0x18, 0x1E, 0x11, 0x19, 0x18, 0x26, 0x5C, 0x00,
	0x58, 0x0E, 0x30, 0x5E, 0x51, 0x25, 0x3C, 0x72, 0x29, 0x2A, 0x22, 0x3E,
	0x01, 0x29, 0x10, 0x1C, 0x03, 0x77, 0x01, 0x0C, 0x1C, 0x1B, 0x2F, 0x0D,
	0x13, 0x59, 0x2C, 0x38, 0x2B, 0x05, 0x28, 0x3D, 0x34, 0x35, 0x14, 0x34,
	0x29, 0x2F, 0x2B, 0x2C, 0x28, 0x5C, 0x21, 0x05, 0x07, 0x3E, 0x23, 0x0E,
	0x0F, 0x0A, 0x04, 0x0F, 0x03, 0x3B, 0x28, 0x5B, 0x06, 0x77, 0x2A, 0x05,
	0x0A, 0x09, 0x37, 0x35, 0x26, 0x08, 0x00, 0x23, 0x55, 0x53, 0x14, 0x38,
	0x30, 0x3D, 0x0F, 0x5A, 0x12, 0x35, 0x2A, 0x54, 0x09, 0x11, 0x33, 0x2A,
	0x50, 0x36, 0x3D, 0x7A, 0x06, 0x34, 0x05, 0x3F, 0x2A, 0x28, 0x32, 0x20,
	0x28, 0x03, 0x1F, 0x15, 0x37, 0x5A, 0x70, 0x1D, 0x11, 0x39, 0x07, 0x0E,
	0x1A, 0x31, 0x2D, 0x33, 0x2E, 0x0B, 0x29, 0x05, 0x5F, 0x13, 0x1A, 0x19,
	0x1A, 0x39, 0x37, 0x05, 0x2F, 0x06, 0x29, 0x06, 0x1C, 0x19, 0x28, 0x24,
	0x10, 0x04, 0x05, 0x3D, 0x04, 0x14, 0x00, 0x05, 0x23, 0x11, 0x00, 0x25,
	0x1B, 0x19, 0x11, 0x77, 0x2B, 0x15, 0x18, 0x1B, 0x6D, 0x1E, 0x05, 0x57,
	0x52, 0x1A, 0x43, 0x0B, 0x28, 0x04, 0x0A, 0x1B, 0x07, 0x3C, 0x5B, 0x36,
	0x36, 0x28, 0x18, 0x04, 0x7B, 0x58, 0x10, 0x41, 0x5D, 0x36, 0x0A, 0x25,
	0x19, 0x27, 0x3A, 0x3A, 0x25, 0x2B, 0x21, 0x0E, 0x47, 0x14, 0x34, 0x0C,
	0x0F, 0x21, 0x2B, 0x5D, 0x33, 0x2E, 0x1D, 0x32, 0x2C, 0x06, 0x13, 0x27,
	0x31, 0x05, 0x27, 0x6D, 0x3D, 0x05, 0x1F, 0x00, 0x6D, 0x2A, 0x55, 0x3C,
	0x52, 0x13, 0x58, 0x33, 0x5B, 0x1E, 0x20, 0x14, 0x07, 0x08, 0x0C, 0x18,
	0x0A, 0x17, 0x26, 0x13, 0x6D, 0x23, 0x56, 0x45, 0x5E, 0x37, 0x35, 0x0A,
	0x2F, 0x31, 0x07, 0x55, 0x0C, 0x22, 0x38, 0x75, 0x5D, 0x3B, 0x37, 0x59,
	0x26, 0x3D, 0x4E, 0x05, 0x3F, 0x30, 0x28, 0x0B, 0x3D, 0x3F, 0x06, 0x1C,
	0x10, 0x17, 0x33, 0x25, 0x3D, 0x53, 0x02, 0x5F, 0x0C, 0x1B, 0x15, 0x22,
	0x2E, 0x76, 0x02, 0x10, 0x1C, 0x5D, 0x38, 0x55, 0x52, 0x18, 0x5C, 0x04,
	0x16, 0x05, 0x0C, 0x3C, 0x16, 0x1A, 0x3B, 0x08, 0x0F, 0x25, 0x0A, 0x2E,
	0x3A, 0x1D, 0x18, 0x3D, 0x0A, 0x28, 0x5A, 0x2B, 0x3E, 0x57, 0x08, 0x24,
	0x26, 0x06, 0x27, 0x34, 0x53, 0x18, 0x01, 0x2B, 0x25, 0x09, 0x18, 0x2F,
	0x27, 0x21, 0x11, 0x21, 0x24, 0x16, 0x3A, 0x3A, 0x11, 0x23, 0x4E, 0x1D,
	0x32, 0x0C, 0x23, 0x09, 0x09, 0x59, 0x73, 0x24, 0x36, 0x14, 0x5C, 0x69,
	0x24, 0x03, 0x0B, 0x44, 0x24, 0x3B, 0x04, 0x45, 0x0C, 0x3B, 0x5F, 0x24,
	0x58, 0x0C, 0x6D, 0x2E, 0x33, 0x00, 0x32, 0x38, 0x1F, 0x25, 0x57, 0x52,
	0x11, 0x5C, 0x4A, 0x3B, 0x01, 0x06, 0x54, 0x2D, 0x5E, 0x1B, 0x7B, 0x36,
	0x31, 0x2A, 0x26, 0x16, 0x2D, 0x0A, 0x5F, 0x5B, 0x36, 0x23, 0x59, 0x18,
	0x12, 0x35, 0x0E, 0x09, 0x21, 0x5F, 0x2B, 0x19, 0x30, 0x1E, 0x5D, 0x7B,
	0x0E, 0x02, 0x0D, 0x1E, 0x6D, 0x5E, 0x51, 0x3E, 0x44, 0x12, 0x55, 0x56,
	0x45, 0x44, 0x27, 0x1E, 0x15, 0x01, 0x5F, 0x15, 0x04, 0x07, 0x5B, 0x0D,
	0x20, 0x2A, 0x29, 0x25, 0x59, 0x21, 0x1E, 0x20, 0x5D, 0x01, 0x1B, 0x2B,
	0x59, 0x1C, 0x20, 0x30, 0x27, 0x32, 0x56, 0x5C, 0x27, 0x3A, 0x54, 0x5C,
	0x3D, 0x1A, 0x02, 0x3B, 0x1D, 0x0D, 0x09, 0x15, 0x10, 0x5B, 0x5D, 0x1A,
	0x34, 0x02, 0x5F, 0x5E, 0x14, 0x0F, 0x12, 0x0C, 0x21, 0x0D, 0x3B, 0x32,
	0x38, 0x5E, 0x2F, 0x28, 0x05, 0x5C, 0x5B, 0x16, 0x39, 0x29, 0x16, 0x5B,
	0x29, 0x0B, 0x53, 0x45, 0x1D, 0x18, 0x5C, 0x2E, 0x0D, 0x1F, 0x1A, 0x2E,
	0x4E, 0x56, 0x53, 0x71, 0x5E, 0x1B, 0x04, 0x5D, 0x03, 0x3A, 0x0A, 0x3B,
	0x28, 0x37, 0x24, 0x29, 0x3A, 0x5F, 0x16, 0x05, 0x22, 0x0B, 0x1C, 0x20,
	0x54, 0x35, 0x2F, 0x13, 0x3B, 0x14, 0x0B, 0x34, 0x5B, 0x77, 0x0D, 0x18,
	0x0C, 0x13, 0x16, 0x05, 0x56, 0x14, 0x29, 0x10, 0x3F, 0x31, 0x0F, 0x18,
	0x2D, 0x23, 0x16, 0x5D, 0x22, 0x00, 0x07, 0x0B, 0x3A, 0x03, 0x29, 0x1D,
	0x16, 0x37, 0x1C, 0x2A, 0x3B, 0x18, 0x0D, 0x25, 0x12, 0x5D, 0x15, 0x02,
	0x04, 0x2F, 0x28, 0x16, 0x2C, 0x5E, 0x1B, 0x1B, 0x50, 0x3B, 0x11, 0x00,
	0x58, 0x26, 0x5E, 0x0C, 0x35, 0x05, 0x14, 0x22, 0x18, 0x32, 0x00, 0x24,
	0x24, 0x3B, 0x36, 0x08, 0x0E, 0x01, 0x19, 0x00, 0x02, 0x57, 0x17, 0x11,
	0x76, 0x06, 0x22, 0x04, 0x2C, 0x0C, 0x1F, 0x28, 0x18, 0x28, 0x32, 0x1C,
	0x2D, 0x39, 0x0E, 0x0B, 0x1A, 0x19, 0x2D, 0x52, 0x38, 0x27, 0x09, 0x23,
	0x03, 0x70, 0x0E, 0x16, 0x04, 0x5E, 0x13, 0x00, 0x24, 0x0C, 0x22, 0x72,
	0x27, 0x24, 0x22, 0x40, 0x20, 0x3F, 0x0F, 0x34, 0x39, 0x28, 0x26, 0x55,
	0x2A, 0x22, 0x09, 0x0B, 0x03, 0x57, 0x5B, 0x74, 0x18, 0x18, 0x2C, 0x22,
	0x69, 0x18, 0x32, 0x1A, 0x53, 0x35, 0x2B, 0x39, 0x3D, 0x5B, 0x14, 0x09,
	0x54, 0x05, 0x29, 0x08, 0x3A, 0x2E, 0x3A, 0x07, 0x06, 0x22, 0x30, 0x07,
	0x3F, 0x2B, 0x01, 0x59, 0x09, 0x08, 0x2E, 0x3B, 0x24, 0x3B, 0x18, 0x07,
	0x00, 0x28, 0x1D, 0x20, 0x2C, 0x09, 0x26, 0x2B, 0x11, 0x07, 0x1D, 0x02,
	0x1D, 0x04, 0x3B, 0x0E, 0x23, 0x01, 0x1C, 0x74, 0x0F, 0x59, 0x1C, 0x3D,
	0x13, 0x20, 0x3B, 0x24, 0x40, 0x06, 0x02, 0x31, 0x3A, 0x2C, 0x11, 0x1D,
	0x38, 0x3E, 0x2A, 0x70, 0x28, 0x51, 0x3F, 0x27, 0x13, 0x04, 0x55, 0x22,
	0x0F, 0x0D, 0x04, 0x31, 0x41, 0x11, 0x29, 0x03, 0x19, 0x3B, 0x21, 0x35,
	0x08, 0x02, 0x45, 0x24, 0x36, 0x3E, 0x13, 0x2B, 0x2E, 0x0B, 0x26, 0x05,
	0x07, 0x1E, 0x70, 0x1B, 0x3B, 0x58, 0x01, 0x01, 0x04, 0x1B, 0x0B, 0x2A,
	0x76, 0x1D, 0x0F, 0x3F, 0x22, 0x17, 0x2B, 0x28, 0x38, 0x20, 0x04, 0x06,
	0x20, 0x01, 0x21, 0x03, 0x04, 0x38, 0x5A, 0x1F, 0x01, 0x2F, 0x55, 0x1F,
	0x0F, 0x06, 0x14, 0x20, 0x5A, 0x20, 0x34, 0x3D, 0x57, 0x37, 0x1D, 0x36,
	0x39, 0x37, 0x26, 0x1D, 0x1B, 0x5B, 0x26, 0x21, 0x02, 0x36, 0x03, 0x11,
	0x19, 0x22, 0x09, 0x27, 0x17, 0x23, 0x5D, 0x01, 0x07, 0x2A, 0x5E, 0x02,
	0x30, 0x14, 0x02, 0x09, 0x5E, 0x09, 0x06, 0x30, 0x1F, 0x3A, 0x21, 0x24,
	0x4E, 0x5F, 0x39, 0x28, 0x5D, 0x51, 0x5B, 0x27, 0x25, 0x2A, 0x28, 0x38,
	0x18, 0x1A, 0x16, 0x06, 0x37, 0x21, 0x29, 0x27, 0x29, 0x3F, 0x00, 0x21,
	0x1E, 0x2A, 0x06, 0x2F, 0x08, 0x14, 0x2F, 0x41, 0x5F, 0x3B, 0x18, 0x2B,
	0x00, 0x2F, 0x08, 0x3A, 0x0F, 0x34, 0x58, 0x75, 0x2D, 0x06, 0x1F, 0x1D,
	0x30, 0x05, 0x0D, 0x00, 0x06, 0x0F, 0x09, 0x2E, 0x5E, 0x3D, 0x07, 0x22,
	0x05, 0x02, 0x1F, 0x26, 0x2E, 0x1B, 0x1F, 0x38, 0x0D, 0x00, 0x2A, 0x5C,
	0x07, 0x20, 0x5C, 0x26, 0x3F, 0x3C, 0x6D, 0x5C, 0x2B, 0x24, 0x33, 0x76,
	0x2D, 0x31, 0x2B, 0x2D, 0x2B, 0x20, 0x52, 0x34, 0x13, 0x29, 0x36, 0x2B,
	0x01, 0x5A, 0x2A, 0x14, 0x2A, 0x2B, 0x22, 0x0C, 0x27, 0x36, 0x45, 0x59,
	0x72, 0x09, 0x0F, 0x1E, 0x08, 0x32, 0x07, 0x04, 0x08, 0x1C, 0x28, 0x1E,
	0x00, 0x04, 0x1B, 0x76, 0x27, 0x57, 0x20, 0x00, 0x76, 0x59, 0x09, 0x5C,
	0x2F, 0x24, 0x0E, 0x28, 0x1A, 0x59, 0x37, 0x39, 0x03, 0x23, 0x12, 0x31,
	0x38, 0x02, 0x0A, 0x59, 0x15, 0x26, 0x37, 0x2C, 0x2C, 0x30, 0x38, 0x2E,
	0x25, 0x1D, 0x28, 0x20, 0x4E, 0x37, 0x0A, 0x1A, 0x1E, 0x00, 0x3C, 0x20,
	0x10, 0x59, 0x52, 0x39, 0x1C, 0x26, 0x55, 0x55, 0x0C, 0x3D, 0x07, 0x18,
	0x13, 0x41, 0x1E, 0x76, 0x2E, 0x09, 0x38, 0x1F, 0x38, 0x20, 0x15, 0x58,
	0x1E, 0x18, 0x05, 0x33, 0x26, 0x11, 0x7B, 0x5C, 0x2B, 0x16, 0x1D, 0x77,
	0x58, 0x04, 0x17, 0x26, 0x16, 0x5F, 0x30, 0x5C, 0x40, 0x00, 0x29, 0x58,
	0x0D, 0x09, 0x3A, 0x0F, 0x56, 0x16, 0x3C, 0x38, 0x2F, 0x22, 0x2A, 0x59,
	0x06, 0x25, 0x37, 0x3D, 0x04, 0x35, 0x0A, 0x33, 0x0B, 0x5E, 0x05, 0x25,
	0x31, 0x3C, 0x1A, 0x16, 0x0D, 0x13, 0x25, 0x39, 0x2C, 0x5D, 0x30, 0x19,
	0x01, 0x1B, 0x28, 0x09, 0x0F, 0x3F, 0x0E, 0x5D, 0x37, 0x0D, 0x1D, 0x76,
	0x5F, 0x23, 0x5B, 0x5B, 0x3B, 0x06, 0x30, 0x38, 0x22, 0x76, 0x01, 0x59,
	0x18, 0x01, 0x16, 0x00, 0x58, 0x0F, 0x3E, 0x12, 0x39, 0x2B, 0x57, 0x19,
	0x0F, 0x5D, 0x2F, 0x5E, 0x39, 0x14, 0x59, 0x24, 0x57, 0x0A, 0x21, 0x3D,
	0x54, 0x3E, 0x33, 0x2E, 0x25, 0x13, 0x0B, 0x3A, 0x07, 0x2A, 0x35, 0x36,
	0x32, 0x24, 0x15, 0x2C, 0x18, 0x38, 0x34, 0x16, 0x02, 0x45, 0x1D, 0x33,
	0x23, 0x0E, 0x17, 0x0D, 0x31, 0x34, 0x05, 0x02, 0x0D, 0x31, 0x0E, 0x31,
	0x19, 0x1E, 0x2A, 0x14, 0x05, 0x0A, 0x20, 0x33, 0x5A, 0x0A, 0x22, 0x06,
	0x18, 0x55, 0x02, 0x0F, 0x38, 0x76, 0x1E, 0x13, 0x19, 0x19, 0x00, 0x0A,
	0x56, 0x36, 0x3C, 0x00, 0x22, 0x1B, 0x0B, 0x06, 0x74, 0x0F, 0x0F, 0x56,
	0x27, 0x09, 0x47, 0x05, 0x06, 0x04, 0x11, 0x54, 0x05, 0x1C, 0x19, 0x2A,
	0x20, 0x16, 0x00, 0x2C, 0x08, 0x0F, 0x38, 0x05, 0x39, 0x2B, 0x34, 0x50,
	0x1F, 0x22, 0x30, 0x00, 0x0B, 0x14, 0x59, 0x34, 0x3A, 0x07, 0x0A, 0x5E,
	0x17, 0x25, 0x35, 0x1C, 0x3A, 0x2D, 0x1A, 0x05, 0x0A, 0x12, 0x1B, 0x2F,
	0x16, 0x57, 0x0F, 0x2B, 0x55, 0x56, 0x04, 0x5E, 0x37, 0x2F, 0x55, 0x5A,
	0x24, 0x2E, 0x1A, 0x34, 0x56, 0x25, 0x27, 0x5E, 0x53, 0x23, 0x13, 0x38,
	0x35, 0x22, 0x01, 0x5E, 0x28, 0x20, 0x0A, 0x58, 0x44, 0x37, 0x25, 0x35,
	0x03, 0x40, 0x29, 0x28, 0x25, 0x27, 0x44, 0x06, 0x16, 0x20, 0x2A, 0x2C,
	0x2A, 0x0F, 0x31, 0x09, 0x05, 0x2B, 0x5F, 0x06, 0x23, 0x2A, 0x10, 0x39,
	0x30, 0x07, 0x38, 0x0A, 0x54, 0x30, 0x24, 0x2C, 0x35, 0x01, 0x27, 0x29,
	0x2A, 0x18, 0x3C, 0x25, 0x37, 0x09, 0x1B, 0x2F, 0x0A, 0x56, 0x0F, 0x2A,
	0x5F, 0x06, 0x28, 0x3F, 0x3B, 0x01, 0x24, 0x0D, 0x25, 0x12, 0x29, 0x52,
	0x18, 0x25, 0x28, 0x21, 0x02, 0x29, 0x2A, 0x33, 0x23, 0x02, 0x16, 0x40,
	0x71, 0x29, 0x19, 0x5E, 0x59, 0x0B, 0x1B, 0x0C, 0x02, 0x21, 0x0E, 0x24,
	0x38, 0x3F, 0x20, 0x00, 0x58, 0x39, 0x21, 0x32, 0x2A, 0x0F, 0x20, 0x27,
	0x24, 0x0F, 0x1B, 0x25, 0x37, 0x28, 0x08, 0x5D, 0x53, 0x28, 0x5C, 0x7B,
	0x2F, 0x0E, 0x17, 0x03, 0x0E, 0x1C, 0x17, 0x3C, 0x03, 0x77, 0x14, 0x05,
	0x58, 0x19, 0x07, 0x36, 0x00, 0x5C, 0x2F, 0x3B, 0x55, 0x2F, 0x03, 0x26,
	0x05, 0x16, 0x20, 0x3D, 0x2A, 0x38, 0x35, 0x0B, 0x5F, 0x26, 0x18, 0x0A,
	0x23, 0x1E, 0x26, 0x38, 0x1F, 0x00, 0x05, 0x1B, 0x1B, 0x1A, 0x18, 0x20,
	0x0C, 0x15, 0x23, 0x03, 0x3D, 0x3D, 0x1B, 0x0A, 0x35, 0x2F, 0x28, 0x26,
	0x07, 0x10, 0x5F, 0x18, 0x08, 0x07, 0x2C, 0x0C, 0x0D, 0x38, 0x55, 0x2D,
	0x26, 0x0C, 0x36, 0x43, 0x26, 0x3A, 0x32, 0x14, 0x09, 0x17, 0x39, 0x28,
	0x16, 0x3B, 0x18, 0x0A, 0x02, 0x26, 0x1E, 0x55, 0x03, 0x58, 0x0A, 0x1F,
	0x34, 0x1F, 0x1C, 0x01, 0x1C, 0x0E, 0x17, 0x3F, 0x7A, 0x01, 0x3B, 0x09,
	0x20, 0x28, 0x0B, 0x57, 0x1C, 0x5F, 0x06, 0x26, 0x2C, 0x39, 0x32, 0x38,
	0x24, 0x00, 0x26, 0x08, 0x2A, 0x0B, 0x51, 0x5A, 0x27, 0x13, 0x2B, 0x38,
	0x3B, 0x0C, 0x74, 0x38, 0x23, 0x2B, 0x13, 0x18, 0x3D, 0x51, 0x58, 0x0F,
	0x1B, 0x1C, 0x50, 0x29, 0x23, 0x09, 0x54, 0x22, 0x27, 0x11, 0x00, 0x04,
	0x2C, 0x56, 0x33, 0x03, 0x58, 0x2B, 0x36, 0x33, 0x33, 0x59, 0x06, 0x14,
	0x24, 0x34, 0x0B, 0x56, 0x0B, 0x2C, 0x38, 0x01, 0x28, 0x37, 0x5E, 0x2E,
	0x15, 0x0C, 0x37, 0x04, 0x7A, 0x28, 0x13, 0x41, 0x2A, 0x75, 0x1F, 0x34,
	0x1B, 0x29, 0x77, 0x58, 0x29, 0x23, 0x32, 0x10, 0x2B, 0x23, 0x23, 0x24,
	0x76, 0x1B, 0x53, 0x23, 0x22, 0x1B, 0x0F, 0x3B, 0x2F, 0x22, 0x35, 0x3A,
	0x09, 0x56, 0x00, 0x03, 0x26, 0x0E, 0x24, 0x00, 0x28, 0x5F, 0x39, 0x3A,
	0x53, 0x08, 0x5C, 0x11, 0x04, 0x18, 0x77, 0x05, 0x39, 0x08, 0x1B, 0x2A,
	0x23, 0x11, 0x0C, 0x24, 0x10, 0x01, 0x20, 0x07, 0x06, 0x75, 0x29, 0x15,
	0x18, 0x2A, 0x77, 0x21, 0x0B, 0x07, 0x3B, 0x08, 0x1D, 0x0C, 0x3B, 0x0F,
	0x05, 0x2A, 0x18, 0x17, 0x06, 0x75, 0x22, 0x50, 0x03, 0x1E, 0x30, 0x04,
	0x50, 0x3F, 0x0D, 0x1B, 0x20, 0x00, 0x2B, 0x0F, 0x0F, 0x22, 0x00, 0x0D,
	0x3C, 0x2C, 0x35, 0x24, 0x1E, 0x1A, 0x11, 0x00, 0x31, 0x2C, 0x09, 0x17,
	0x21, 0x0F, 0x58, 0x53, 0x05, 0x01, 0x39, 0x14, 0x59, 0x0D, 0x02, 0x55,
	0x09, 0x5B, 0x74, 0x36, 0x26, 0x34, 0x18, 0x08, 0x1B, 0x52, 0x03, 0x31,
	0x31, 0x59, 0x0C, 0x06, 0x3C, 0x09, 0x0F, 0x37, 0x03, 0x5E, 0x29, 0x2D,
	0x35, 0x29, 0x39, 0x30, 0x08, 0x14, 0x5A, 0x19, 0x25, 0x0F, 0x0C, 0x16,
	0x32, 0x0D, 0x1F, 0x02, 0x2C, 0x28, 0x23, 0x3C, 0x16, 0x5B, 0x1C, 0x06,
	0x3E, 0x0C, 0x2A, 0x21, 0x28, 0x1A, 0x34, 0x37, 0x2C, 0x00, 0x47, 0x2E,
	0x08, 0x52, 0x11, 0x0B, 0x23, 0x5F, 0x38, 0x70, 0x35, 0x04, 0x1D, 0x32,
	0x1B, 0x1F, 0x00, 0x39, 0x11, 0x18, 0x0B, 0x23, 0x5E, 0x5E, 0x32, 0x38,
	0x34, 0x07, 0x0F, 0x25, 0x09, 0x23, 0x14, 0x2C, 0x03, 0x59, 0x06, 0x25,
	0x3F, 0x2E, 0x1F, 0x2F, 0x2C, 0x2A, 0x1B, 0x43, 0x14, 0x17, 0x39, 0x0E,
	0x26, 0x16, 0x0F, 0x44, 0x0C, 0x5E, 0x0B, 0x0C, 0x04, 0x1B, 0x21, 0x2D,
	0x24, 0x44, 0x21, 0x35, 0x51, 0x21, 0x05, 0x05, 0x35, 0x38, 0x0C, 0x3E,
	0x2D, 0x14, 0x58, 0x5C, 0x31, 0x0C, 0x34, 0x39, 0x29, 0x2C, 0x01, 0x0F,
	0x2E, 0x2A, 0x19, 0x16, 0x0B, 0x02, 0x03, 0x59, 0x18, 0x5D, 0x14, 0x5A,
	0x29, 0x00, 0x05, 0x39, 0x3A, 0x06, 0x3A, 0x01, 0x20, 0x14, 0x2A, 0x69,
	0x24, 0x20, 0x18, 0x44, 0x3A, 0x06, 0x38, 0x59, 0x18, 0x2C, 0x34, 0x2E,
	0x2F, 0x21, 0x12, 0x02, 0x19, 0x29, 0x31, 0x37, 0x58, 0x0D, 0x25, 0x53,
	0x18, 0x54, 0x05, 0x58, 0x01, 0x20, 0x5F, 0x33, 0x04, 0x3F, 0x0C, 0x19,
	0x16, 0x2F, 0x03, 0x10, 0x5E, 0x3B, 0x5D, 0x25, 0x7A, 0x25, 0x27, 0x2C,
	0x3B, 0x26, 0x05, 0x2C, 0x25, 0x11, 0x00, 0x3B, 0x0F, 0x20, 0x12, 0x28,
	0x0B, 0x32, 0x00, 0x19, 0x3B, 0x08, 0x03, 0x24, 0x2A, 0x33, 0x0D, 0x34,
	0x5A, 0x5C, 0x0A, 0x1C, 0x16, 0x21, 0x11, 0x25, 0x14, 0x27, 0x01, 0x2E,
	0x28, 0x21, 0x22, 0x38, 0x33, 0x23, 0x0A, 0x29, 0x0D, 0x2D, 0x77, 0x19,
	0x29, 0x24, 0x1E, 0x00, 0x15, 0x39, 0x34, 0x05, 0x0F, 0x5C, 0x4A, 0x2C,
	0x20, 0x24, 0x2A, 0x0F, 0x23, 0x13, 0x69, 0x2E, 0x18, 0x3F, 0x1F, 0x2A,
	0x21, 0x52, 0x01, 0x1C, 0x33, 0x07, 0x0A, 0x5A, 0x0E, 0x20, 0x39, 0x27,
	0x24, 0x04, 0x2C, 0x28, 0x05, 0x2F, 0x3D, 0x05, 0x1B, 0x26, 0x2B, 0x28,
	0x25, 0x25, 0x0F, 0x09, 0x26, 0x01, 0x26, 0x06, 0x2B, 0x01, 0x25, 0x21,
	0x39, 0x04, 0x01, 0x3A, 0x2B, 0x59, 0x0B, 0x23, 0x76, 0x58, 0x22, 0x24,
	0x5E, 0x0D, 0x0B, 0x12, 0x2F, 0x40, 0x1B, 0x08, 0x33, 0x5C, 0x08, 0x06,
	0x21, 0x28, 0x1D, 0x5F, 0x24, 0x0A, 0x20, 0x5A, 0x26, 0x12, 0x14, 0x23,
	0x59, 0x27, 0x0B, 0x43, 0x20, 0x58, 0x32, 0x29, 0x05, 0x37, 0x5C, 0x20,
	0x75, 0x59, 0x09, 0x24, 0x31, 0x37, 0x19, 0x51, 0x09, 0x27, 0x05, 0x36,
	0x0D, 0x56, 0x21, 0x2F, 0x3C, 0x28, 0x26, 0x21, 0x16, 0x01, 0x39, 0x26,
	0x2E, 0x37, 0x2E, 0x2B, 0x2D, 0x53, 0x24, 0x16, 0x20, 0x5A, 0x2F, 0x2A,
	0x1C, 0x56, 0x28, 0x5A, 0x29, 0x03, 0x20, 0x16, 0x3F, 0x05, 0x0F, 0x1B,
	0x27, 0x5F, 0x07, 0x1C, 0x54, 0x24, 0x39, 0x2B, 0x26, 0x0A, 0x58, 0x31,
	0x35, 0x15, 0x16, 0x29, 0x1B, 0x32, 0x26, 0x35, 0x1C, 0x05, 0x3A, 0x0B,
	0x32, 0x04, 0x00, 0x74, 0x3B, 0x55, 0x2A, 0x31, 0x2D, 0x5E, 0x25, 0x07,
	0x26, 0x38, 0x22, 0x27, 0x45, 0x2E, 0x15, 0x01, 0x22, 0x01, 0x5C, 0x0D,
	0x0A, 0x15, 0x2C, 0x5E, 0x38, 0x07, 0x0F, 0x00, 0x2C, 0x28, 0x2F, 0x31,
	0x21, 0x3A, 0x38, 0x47, 0x27, 0x09, 0x01, 0x69, 0x04, 0x0A, 0x2C, 0x3D,
	0x11, 0x0A, 0x24, 0x25, 0x1C, 0x08, 0x54, 0x55, 0x21, 0x1E, 0x70, 0x22,
	0x59, 0x22, 0x08, 0x14, 0x5E, 0x2D, 0x5D, 0x21, 0x01, 0x36, 0x08, 0x25,
	0x09, 0x0B, 0x58, 0x52, 0x09, 0x23, 0x07, 0x36, 0x1B, 0x5E, 0x5E, 0x0A,
	0x0B, 0x09, 0x03, 0x24, 0x12, 0x08, 0x0F, 0x2F, 0x24, 0x0A, 0x2B, 0x38,
	0x1B, 0x08, 0x06, 0x1B, 0x2E, 0x0D, 0x1C, 0x33, 0x35, 0x2F, 0x2C, 0x3E,
	0x26, 0x1F, 0x13, 0x0C, 0x0C, 0x0F, 0x02, 0x0B, 0x00, 0x24, 0x0F, 0x23,
	0x20, 0x02, 0x3B, 0x09, 0x35, 0x34, 0x5A, 0x2F, 0x29, 0x16, 0x2E, 0x26,
	0x26, 0x71, 0x21, 0x20, 0x5B, 0x03, 0x11, 0x02, 0x05, 0x00, 0x3F, 0x25,
	0x06, 0x2A, 0x08, 0x2D, 0x05, 0x3D, 0x26, 0x0F, 0x2A, 0x3A, 0x23, 0x3B,
	0x17, 0x5F, 0x75, 0x00, 0x22, 0x01, 0x13, 0x25, 0x3C, 0x11, 0x1B, 0x21,
	0x00, 0x5A, 0x3B, 0x07, 0x22, 0x15, 0x08, 0x02, 0x2C, 0x38, 0x23, 0x24,
	0x0A, 0x41, 0x18, 0x29, 0x1E, 0x27, 0x3E, 0x2A, 0x73, 0x00, 0x0A, 0x22,
	0x3F, 0x04, 0x58, 0x2B, 0x34, 0x5B, 0x76, 0x2F, 0x35, 0x23, 0x00, 0x2F,
	0x08, 0x13, 0x00, 0x24, 0x76, 0x1E, 0x16, 0x5C, 0x18, 0x71, 0x34, 0x16,
	0x5A, 0x1A, 0x0A, 0x36, 0x36, 0x57, 0x01, 0x0F, 0x26, 0x53, 0x2A, 0x5F,
	0x10, 0x16, 0x08, 0x5F, 0x2A, 0x70, 0x08, 0x11, 0x02, 0x5C, 0x0C, 0x1F,
	0x19, 0x09, 0x5F, 0x1B, 0x5F, 0x0B, 0x05, 0x59, 0x76, 0x1B, 0x57, 0x23,
	0x5F, 0x09, 0x20, 0x18, 0x3E, 0x2D, 0x35, 0x5E, 0x10, 0x58, 0x3F, 0x2C,
	0x58, 0x33, 0x2D, 0x0D, 0x37, 0x5C, 0x32, 0x2B, 0x0D, 0x00, 0x5B, 0x2E,
	0x3F, 0x44, 0x08, 0x59, 0x2E, 0x2A, 0x5C, 0x20, 0x39, 0x38, 0x07, 0x01,
	0x35, 0x54, 0x1B, 0x2A, 0x53, 0x77, 0x2E, 0x59, 0x26, 0x07, 0x75, 0x15,
	0x0F, 0x05, 0x3F, 0x21, 0x38, 0x35, 0x5A, 0x3B, 0x3A, 0x43, 0x05, 0x0D,
	0x31, 0x12, 0x3C, 0x16, 0x5D, 0x2C, 0x2D, 0x34, 0x38, 0x3E, 0x21, 0x77,
	0x23, 0x2D, 0x5B, 0x58, 0x0B, 0x59, 0x14, 0x26, 0x0E, 0x74, 0x06, 0x09,
	0x20, 0x39, 0x72, 0x58, 0x2E, 0x1D, 0x1C, 0x7A, 0x34, 0x28, 0x2A, 0x00,
	0x21, 0x5E, 0x18, 0x1C, 0x40, 0x30, 0x27, 0x13, 0x22, 0x24, 0x76, 0x3B,
	0x38, 0x3D, 0x1C, 0x6D, 0x59, 0x53, 0x25, 0x0F, 0x00, 0x18, 0x36, 0x21,
	0x5F, 0x3B, 0x5C, 0x04, 0x0A, 0x3B, 0x33, 0x1E, 0x18, 0x45, 0x58, 0x3A,
	0x1D, 0x27, 0x2B, 0x05, 0x72, 0x5D, 0x06, 0x5C, 0x2C, 0x77, 0x0E, 0x3B,
	0x37, 0x5F, 0x0E, 0x07, 0x05, 0x14, 0x05, 0x1B, 0x2B, 0x54, 0x59, 0x11,
	0x10, 0x55, 0x38, 0x16, 0x5E, 0x77, 0x0A, 0x31, 0x56, 0x2E, 0x27, 0x1E,
	0x0C, 0x21, 0x23, 0x6D, 0x05, 0x04, 0x18, 0x19, 0x11, 0x18, 0x51, 0x14,
	0x44, 0x08, 0x3B, 0x55, 0x36, 0x2D, 0x24, 0x35, 0x13, 0x39, 0x3E, 0x24,
	0x1E, 0x17, 0x0A, 0x12, 0x0C, 0x02, 0x2C, 0x20, 0x06, 0x07, 0x03, 0x2E,
	0x56, 0x1C, 0x05, 0x35, 0x17, 0x25, 0x1F, 0x31, 0x1C, 0x06, 0x03, 0x5F,
	0x32, 0x25, 0x35, 0x2A, 0x0F, 0x03, 0x0D, 0x0C, 0x02, 0x26, 0x0D, 0x58,
	0x20, 0x5F, 0x3B, 0x05, 0x35, 0x34, 0x25, 0x29, 0x33, 0x09, 0x30, 0x19,
	0x0C, 0x76, 0x28, 0x2B, 0x18, 0x18, 0x18, 0x01, 0x59, 0x3E, 0x0E, 0x00,
	0x3F, 0x0B, 0x00, 0x26, 0x03, 0x1C, 0x1B, 0x36, 0x39, 0x71, 0x0D, 0x4E,
	0x39, 0x22, 0x26, 0x38, 0x17, 0x1D, 0x31, 0x37, 0x01, 0x39, 0x56, 0x2F,
	0x35, 0x5B, 0x17, 0x21, 0x01, 0x2C, 0x39, 0x25, 0x1E, 0x53, 0x3A, 0x04,
	0x15, 0x3E, 0x2A, 0x3B, 0x19, 0x02, 0x5E, 0x32, 0x12, 0x55, 0x2F, 0x23,
	0x2C, 0x70, 0x2E, 0x55, 0x28, 0x31, 0x38, 0x3E, 0x23, 0x06, 0x02, 0x1A,
	0x1C, 0x0C, 0x19, 0x0F, 0x07, 0x38, 0x25, 0x5A, 0x3C, 0x38, 0x5D, 0x37,
	0x3A, 0x2F, 0x0B, 0x1B, 0x54, 0x0F, 0x31, 0x31, 0x36, 0x08, 0x14, 0x3C,
	0x76, 0x38, 0x23, 0x14, 0x08, 0x16, 0x03, 0x02, 0x24, 0x03, 0x6D, 0x1E,
	0x02, 0x28, 0x27, 0x27, 0x2E, 0x0A, 0x19, 0x2D, 0x1A, 0x1D, 0x27, 0x36,
	0x3E, 0x1B, 0x03, 0x35, 0x21, 0x29, 0x20, 0x2A, 0x3B, 0x07, 0x5E, 0x2B,
	0x01, 0x59, 0x3E, 0x00, 0x20, 0x0D, 0x2E, 0x39, 0x40, 0x38, 0x0D, 0x06,
	0x2B, 0x13, 0x2E, 0x09, 0x15, 0x5E, 0x5F, 0x06, 0x01, 0x25, 0x1A, 0x33,
	0x2A, 0x18, 0x00, 0x1A, 0x5B, 0x35, 0x5D, 0x51, 0x0D, 0x07, 0x16, 0x07,
	0x2B, 0x3F, 0x0A, 0x26, 0x29, 0x09, 0x36, 0x58, 0x2D, 0x5A, 0x00, 0x2D,
	0x3F, 0x32, 0x58, 0x2A, 0x00, 0x0E, 0x70, 0x0B, 0x16, 0x57, 0x26, 0x25,
	0x3B, 0x2B, 0x58, 0x44, 0x25, 0x24, 0x31, 0x36, 0x07, 0x08, 0x08, 0x58,
	0x25, 0x3B, 0x12, 0x15, 0x12, 0x2B, 0x28, 0x0A, 0x5B, 0x38, 0x5E, 0x5C,
	0x2D, 0x2A, 0x2E, 0x06, 0x13, 0x70, 0x35, 0x10, 0x09, 0x0E, 0x07, 0x0E,
	0x12, 0x24, 0x07, 0x74, 0x06, 0x34, 0x26, 0x23, 0x25, 0x26, 0x50, 0x17,
	0x21, 0x70, 0x2D, 0x04, 0x0D, 0x53, 0x20, 0x02, 0x20, 0x25, 0x11, 0x06,
	0x35, 0x36, 0x25, 0x29, 0x3B, 0x38, 0x27, 0x05, 0x1B, 0x38, 0x21, 0x22,
	0x29, 0x26, 0x12, 0x5A, 0x56, 0x26, 0x3A, 0x2F, 0x22, 0x59, 0x34, 0x33,
	0x07, 0x5E, 0x18, 0x0A, 0x13, 0x1B, 0x5F, 0x19, 0x5F, 0x32, 0x10, 0x0F,
	0x33, 0x14, 0x3A, 0x17, 0x1A, 0x1B, 0x3D, 0x24, 0x14, 0x1B, 0x0D, 0x04,
	0x13, 0x3B, 0x1E, 0x22, 0x1D, 0x3D, 0x16, 0x0F, 0x0F, 0x0C, 0x1E, 0x0D,
	0x0F, 0x50, 0x0B, 0x03, 0x2D, 0x58, 0x02, 0x26, 0x2F, 0x72, 0x58, 0x17,
	0x0F, 0x2A, 0x36, 0x21, 0x08, 0x37, 0x1B, 0x1B, 0x25, 0x00, 0x2A, 0x2F,
	0x17, 0x5D, 0x24, 0x36, 0x2E, 0x71, 0x28, 0x2A, 0x25, 0x05, 0x13, 0x5E,
	0x06, 0x05, 0x5D, 0x04, 0x05, 0x13, 0x14, 0x1E, 0x25, 0x03, 0x57, 0x06,
	0x02, 0x2C, 0x3D, 0x2C, 0x56, 0x29, 0x27, 0x15, 0x37, 0x25, 0x38, 0x06,
	0x1A, 0x56, 0x2D, 0x3D, 0x3A, 0x15, 0x0C, 0x1E, 0x2E, 0x0F, 0x0A, 0x08,
	0x5F, 0x25, 0x26, 0x0B, 0x38, 0x26, 0x0C, 0x21, 0x02, 0x38, 0x00, 0x2A,
	0x10, 0x24, 0x2A, 0x37, 0x1E, 0x21, 0x2E, 0x0A, 0x0D, 0x53, 0x21, 0x22,
	0x38, 0x26, 0x22, 0x76, 0x16, 0x20, 0x5B, 0x0C, 0x69, 0x2E, 0x1B, 0x03,
	0x27, 0x06, 0x2D, 0x22, 0x2A, 0x1D, 0x0F, 0x3D, 0x26, 0x2C, 0x08, 0x0D,
	0x54, 0x19, 0x39, 0x05, 0x0B, 0x5E, 0x2A, 0x5D, 0x29, 0x03, 0x5F, 0x0E,
	0x5C, 0x38, 0x17, 0x0F, 0x11, 0x07, 0x26, 0x35, 0x07, 0x08, 0x36, 0x18,
	0x2E, 0x18, 0x22, 0x04, 0x20, 0x23, 0x27, 0x4E, 0x18, 0x07, 0x17, 0x5D,
	0x20, 0x01, 0x3A, 0x03, 0x0B, 0x19, 0x3C, 0x26, 0x08, 0x1A, 0x56, 0x34,
	0x2A, 0x74, 0x3F, 0x02, 0x1C, 0x0E, 0x3A, 0x5C, 0x55, 0x05, 0x2A, 0x2C,
	0x3E, 0x51, 0x36, 0x1D, 0x38, 0x0B, 0x36, 0x0A, 0x38, 0x2A, 0x39, 0x58,
	0x28, 0x5F, 0x7A, 0x55, 0x2E, 0x36, 0x33, 0x17, 0x06, 0x17, 0x16, 0x18,
	0x0E, 0x06, 0x14, 0x2A, 0x32, 0x08, 0x5E, 0x2F, 0x1A, 0x13, 0x06, 0x5A,
	0x13, 0x27, 0x5E, 0x1B, 0x01, 0x4E, 0x16, 0x18, 0x2C, 0x05, 0x53, 0x08,
	0x18, 0x3A, 0x29, 0x33, 0x2A, 0x31, 0x0A, 0x3F, 0x2B, 0x04, 0x40, 0x20,
	0x3E, 0x59, 0x1C, 0x19, 0x2B, 0x1B, 0x08, 0x1E, 0x0F, 0x2B, 0x5A, 0x32,
	0x00, 0x53, 0x71, 0x16, 0x27, 0x29, 0x0D, 0x12, 0x08, 0x58, 0x38, 0x5A,
	0x2F, 0x20, 0x2E, 0x5B, 0x06, 0x30, 0x1E, 0x59, 0x59, 0x21, 0x29, 0x22,
	0x2E, 0x1E, 0x2D, 0x21, 0x24, 0x04, 0x34, 0x18, 0x2C, 0x00, 0x50, 0x08,
	0x33, 0x33, 0x58, 0x28, 0x34, 0x11, 0x2B, 0x28, 0x2A, 0x2D, 0x0F, 0x04,
	0x02, 0x53, 0x28, 0x27, 0x24, 0x19, 0x24, 0x23, 0x40, 0x72, 0x34, 0x27,
	0x29, 0x3D, 0x1B, 0x38, 0x33, 0x18, 0x3A, 0x09, 0x1C, 0x0F, 0x34, 0x1A,
	0x0D, 0x54, 0x2F, 0x0F, 0x0C, 0x2D, 0x59, 0x24, 0x3C, 0x33, 0x71, 0x5D,
	0x23, 0x1E, 0x5B, 0x11, 0x2A, 0x07, 0x3B, 0x5A, 0x0A, 0x02, 0x32, 0x17,
	0x3D, 0x23, 0x3F, 0x1B, 0x26, 0x05, 0x10, 0x27, 0x37, 0x0F, 0x39, 0x38,
	0x2F, 0x52, 0x3A, 0x12, 0x36, 0x1E, 0x29, 0x0C, 0x5F, 0x17, 0x08, 0x12,
	0x01, 0x32, 0x32, 0x35, 0x23, 0x00, 0x28, 0x27, 0x16, 0x27, 0x21, 0x39,
	0x37, 0x1B, 0x52, 0x39, 0x59, 0x21, 0x2A, 0x2E, 0x1B, 0x39, 0x26, 0x01,
	0x37, 0x25, 0x3A, 0x31, 0x2E, 0x33, 0x5F, 0x2F, 0x04, 0x38, 0x10, 0x1C,
	0x3A, 0x01, 0x08, 0x32, 0x06, 0x08, 0x76, 0x1C, 0x51, 0x2C, 0x23, 0x17,
	0x03, 0x32, 0x21, 0x5C, 0x2D, 0x19, 0x4A, 0x27, 0x21, 0x2C, 0x14, 0x08,
	0x57, 0x52, 0x38, 0x24, 0x24, 0x29, 0x18, 0x11, 0x04, 0x58, 0x28, 0x18,
	0x28, 0x1A, 0x20, 0x2D, 0x26, 0x1A, 0x34, 0x0C, 0x5F, 0x3A, 0x0C, 0x5C,
	0x18, 0x02, 0x3F, 0x1B, 0x29, 0x16, 0x56, 0x5D, 0x24, 0x2E, 0x39, 0x1E,
	0x11, 0x0F, 0x3E, 0x54, 0x1F, 0x0D, 0x25, 0x08, 0x3B, 0x2F, 0x44, 0x2D,
	0x19, 0x2A, 0x04, 0x22, 0x74, 0x16, 0x56, 0x01, 0x31, 0x00, 0x55, 0x06,
	0x0B, 0x5A, 0x76, 0x3C, 0x33, 0x06, 0x2D, 0x06, 0x2A, 0x03, 0x05, 0x5C,
	0x25, 0x39, 0x57, 0x5C, 0x1A, 0x2E, 0x27, 0x20, 0x04, 0x00, 0x00, 0x2A,
	0x2E, 0x1B, 0x24, 0x3A, 0x16, 0x0A, 0x28, 0x59, 0x75, 0x1D, 0x14, 0x2C,
	0x00, 0x10, 0x14, 0x0C, 0x04, 0x5A, 0x33, 0x5B, 0x06, 0x2D, 0x00, 0x75,
	0x1B, 0x0C, 0x34, 0x1E, 0x03, 0x47, 0x2F, 0x17, 0x01, 0x0F, 0x5E, 0x59,
	0x2F, 0x5D, 0x20, 0x05, 0x2E, 0x21, 0x0D, 0x21, 0x5F, 0x33, 0x24, 0x53,
	0x33, 0x21, 0x2D, 0x2D, 0x25, 0x2E, 0x06, 0x0F, 0x24, 0x2F, 0x37, 0x3B,
	0x26, 0x14, 0x2A, 0x14, 0x1C, 0x58, 0x03, 0x26, 0x01, 0x26, 0x09, 0x25,
	0x2D, 0x23, 0x3B, 0x38, 0x5D, 0x39, 0x08, 0x0A, 0x56, 0x59, 0x29, 0x28,
	0x0E, 0x30, 0x2F, 0x06, 0x30, 0x58, 0x1B, 0x20, 0x23, 0x0F, 0x0F, 0x11,
	0x1F, 0x5C, 0x01, 0x02, 0x24, 0x00, 0x39, 0x09, 0x3A, 0x2E, 0x3A, 0x3D,
	0x2F, 0x2D, 0x05, 0x5B, 0x33, 0x15, 0x27, 0x0F, 0x0C, 0x2A, 0x70, 0x21,
	0x06, 0x23, 0x25, 0x07, 0x2D, 0x2C, 0x20, 0x3F, 0x29, 0x08, 0x05, 0x37,
	0x5B, 0x01, 0x07, 0x13, 0x5B, 0x53, 0x3A, 0x2D, 0x2C, 0x26, 0x24, 0x14,
	0x16, 0x04, 0x19, 0x2E, 0x32, 0x19, 0x30, 0x0F, 0x06, 0x75, 0x07, 0x22,
	0x3A, 0x21, 0x74, 0x27, 0x02, 0x45, 0x5F, 0x75, 0x5C, 0x28, 0x03, 0x53,
	0x3B, 0x35, 0x54, 0x38, 0x58, 0x35, 0x14, 0x32, 0x38, 0x03, 0x05, 0x1E,
	0x2E, 0x45, 0x01, 0x29, 0x5F, 0x26, 0x08, 0x23, 0x01, 0x0B, 0x00, 0x03,
	0x53, 0x25, 0x2B, 0x03, 0x3D, 0x3A, 0x09, 0x01, 0x37, 0x2B, 0x3E, 0x74,
	0x0F, 0x59, 0x5C, 0x1C, 0x0B, 0x16, 0x0C, 0x02, 0x2A, 0x0B, 0x0D, 0x17,
	0x37, 0x02, 0x75, 0x14, 0x23, 0x25, 0x0D, 0x7A, 0x04, 0x09, 0x5C, 0x27,
	0x0F, 0x03, 0x04, 0x17, 0x0D, 0x70, 0x25, 0x1B, 0x02, 0x18, 0x00, 0x07,
	0x07, 0x5C, 0x08, 0x38, 0x5F, 0x38, 0x2B, 0x1B, 0x69, 0x54, 0x0D, 0x03,
	0x2A, 0x31, 0x16, 0x19, 0x38, 0x11, 0x36, 0x26, 0x27, 0x04, 0x26, 0x03,
	0x2B, 0x23, 0x59, 0x21, 0x18, 0x18, 0x2A, 0x2F, 0x00, 0x23, 0x05, 0x1B,
	0x03, 0x39, 0x3A, 0x0B, 0x39, 0x3E, 0x3F, 0x1B, 0x16, 0x23, 0x1E, 0x0C,
	0x00, 0x3C, 0x39, 0x37, 0x11, 0x06, 0x59, 0x06, 0x3D, 0x07, 0x15, 0x5C,
	0x0B, 0x36, 0x1D, 0x1B, 0x24, 0x09, 0x3B, 0x5D, 0x15, 0x1D, 0x53, 0x09,
	0x23, 0x23, 0x1E, 0x30, 0x0F, 0x3A, 0x31, 0x5A, 0x2D, 0x07, 0x1B, 0x72,
	0x3D, 0x0A, 0x2D, 0x23, 0x32, 0x5C, 0x2B, 0x00, 0x2F, 0x0D, 0x0B, 0x06,
	0x37, 0x58, 0x1B, 0x1C, 0x54, 0x09, 0x25, 0x16, 0x15, 0x11, 0x00, 0x44,
	0x04, 0x2D, 0x2A, 0x3A, 0x19, 0x10, 0x04, 0x27, 0x5B, 0x3F, 0x0F, 0x24,
	0x53, 0x34, 0x00, 0x10, 0x1C, 0x56, 0x16, 0x2D, 0x00, 0x2A, 0x04, 0x0F,
	0x05, 0x12, 0x23, 0x0B, 0x08, 0x24, 0x18, 0x3D, 0x51, 0x38, 0x0C, 0x69,
	0x0F, 0x51, 0x2A, 0x3D, 0x0C, 0x1A, 0x0F, 0x23, 0x3A, 0x18, 0x29, 0x39,
	0x0D, 0x0A, 0x33, 0x5A, 0x25, 0x04, 0x25, 0x38, 0x15, 0x2F, 0x38, 0x3E,
	0x1A, 0x24, 0x02, 0x1C, 0x58, 0x3B, 0x1C, 0x30, 0x14, 0x29, 0x35, 0x01,
	0x00, 0x25, 0x02, 0x27, 0x23, 0x37, 0x3A, 0x5F, 0x3B, 0x5B, 0x50, 0x3C,
	0x04, 0x23, 0x5A, 0x02, 0x2A, 0x1F, 0x75, 0x1B, 0x1B, 0x2F, 0x2C, 0x6D,
	0x38, 0x0D, 0x1C, 0x19, 0x38, 0x25, 0x24, 0x1E, 0x0E, 0x73, 0x59, 0x25,
	0x5B, 0x07, 0x77, 0x2E, 0x58, 0x34, 0x21, 0x15, 0x5F, 0x05, 0x45, 0x04,
	0x7A, 0x00, 0x06, 0x07, 0x3D, 0x2F, 0x1E, 0x15, 0x21, 0x20, 0x3B, 0x14,
	0x56, 0x28, 0x0F, 0x27, 0x2E, 0x05, 0x21, 0x1B, 0x2F, 0x58, 0x38, 0x3D,
	0x5F, 0x3A, 0x2F, 0x2D, 0x02, 0x21, 0x28, 0x23, 0x25, 0x08, 0x3A, 0x17,
	0x28, 0x25, 0x20, 0x1D, 0x72, 0x3F, 0x2D, 0x02, 0x53, 0x77, 0x0D, 0x55,
	0x1F, 0x26, 0x04, 0x05, 0x13, 0x01, 0x3E, 0x08, 0x1F, 0x0E, 0x39, 0x08,
	0x17, 0x2A, 0x34, 0x58, 0x08, 0x26, 0x27, 0x24, 0x04, 0x21, 0x16, 0x2E,
	0x02, 0x22, 0x5A, 0x1A, 0x00, 0x33, 0x0A, 0x3F, 0x2B, 0x04, 0x2B, 0x5B,
	0x20, 0x15, 0x1D, 0x10, 0x00, 0x33, 0x7B, 0x3D, 0x06, 0x5A, 0x1A, 0x11,
	0x5D, 0x10, 0x3F, 0x01, 0x09, 0x1B, 0x39, 0x57, 0x5A, 0x28, 0x2F, 0x05,
	0x21, 0x58, 0x73, 0x5F, 0x09, 0x0F, 0x1B, 0x08, 0x1C, 0x52, 0x1C, 0x31,
	0x70, 0x0A, 0x54, 0x06, 0x12, 0x36, 0x5A, 0x0E, 0x04, 0x19, 0x0E, 0x43,
	0x27, 0x56, 0x19, 0x2E, 0x07, 0x2A, 0x3F, 0x04, 0x14, 0x1B, 0x53, 0x41,
	0x24, 0x06, 0x23, 0x0D, 0x56, 0x25, 0x00, 0x3D, 0x10, 0x0B, 0x26, 0x76,
	0x39, 0x15, 0x5A, 0x59, 0x2B, 0x24, 0x13, 0x38, 0x0F, 0x18, 0x05, 0x18,
	0x39, 0x12, 0x34, 0x27, 0x29, 0x06, 0x53, 0x16, 0x0B, 0x57, 0x56, 0x0E,
	0x2E, 0x2E, 0x55, 0x23, 0x59, 0x7B, 0x22, 0x2A, 0x36, 0x05, 0x18, 0x09,
	0x0B, 0x0C, 0x40, 0x36, 0x3F, 0x54, 0x09, 0x3B, 0x29, 0x2A, 0x04, 0x5F,
	0x3D, 0x20, 0x15, 0x05, 0x09, 0x3D, 0x2B, 0x1A, 0x26, 0x1C, 0x21, 0x0A,
	0x0B, 0x20, 0x1E, 0x0C, 0x69, 0x2F, 0x13, 0x03, 0x27, 0x26, 0x55, 0x03,
	0x1D, 0x3D, 0x37, 0x58, 0x32, 0x2D, 0x38, 0x75, 0x01, 0x28, 0x02, 0x1D,
	0x08, 0x29, 0x4A, 0x00, 0x0E, 0x2E, 0x5F, 0x02, 0x3C, 0x1F, 0x15, 0x09,
	0x36, 0x25, 0x03, 0x15, 0x2A, 0x1B, 0x3B, 0x53, 0x69, 0x3A, 0x22, 0x1A,
	0x27, 0x2F, 0x1C, 0x55, 0x2B, 0x04, 0x0F, 0x36, 0x2B, 0x0D, 0x1A, 0x73,
	0x3A, 0x07, 0x57, 0x1A, 0x30, 0x5A, 0x38, 0x02, 0x23, 0x3B, 0x3B, 0x16,
	0x3A, 0x1D, 0x17, 0x5B, 0x06, 0x36, 0x0C, 0x07, 0x29, 0x2F, 0x3F, 0x5A,
	0x03, 0x06, 0x23, 0x5F, 0x5B, 0x14, 0x00, 0x33, 0x28, 0x12, 0x2E, 0x3E,
	0x34, 0x18, 0x1B, 0x08, 0x1C, 0x57, 0x1C, 0x20, 0x29, 0x26, 0x02, 0x57,
	0x1B, 0x77, 0x24, 0x10, 0x0A, 0x07, 0x28, 0x26, 0x2A, 0x0C, 0x1E, 0x11,
	0x28, 0x0D, 0x3E, 0x59, 0x29, 0x06, 0x13, 0x0F, 0x04, 0x26, 0x16, 0x0C,
	0x18, 0x2D, 0x69, 0x1B, 0x53, 0x3B, 0x3D, 0x2A, 0x0F, 0x53, 0x34, 0x02,
	0x17, 0x01, 0x19, 0x23, 0x3D, 0x04, 0x1E, 0x12, 0x08, 0x59, 0x1B, 0x16,
	0x07, 0x00, 0x39, 0x12, 0x36, 0x0F, 0x3E, 0x1F, 0x16, 0x54, 0x39, 0x56,
	0x02, 0x31, 0x5E, 0x37, 0x18, 0x59, 0x00, 0x16, 0x2D, 0x5A, 0x33, 0x0C,
	0x09, 0x2A, 0x5E, 0x53, 0x34, 0x2A, 0x35, 0x0B, 0x0D, 0x70, 0x0D, 0x1B,
	0x01, 0x32, 0x2C, 0x1D, 0x4E, 0x02, 0x5E, 0x11, 0x3E, 0x19, 0x1B, 0x3F,
	0x70, 0x47, 0x16, 0x17, 0x3A, 0x0E, 0x34, 0x2F, 0x0F, 0x3A, 0x33, 0x0E,
	0x11, 0x3B, 0x05, 0x32, 0x5A, 0x33, 0x05, 0x38, 0x26, 0x06, 0x02, 0x38,
	0x02, 0x1B, 0x0E, 0x27, 0x07, 0x1A, 0x08, 0x07, 0x05, 0x58, 0x3F, 0x32,
	0x1C, 0x52, 0x5F, 0x00, 0x38, 0x24, 0x25, 0x34, 0x2E, 0x6D, 0x0F, 0x18,
	0x2C, 0x06, 0x6D, 0x0D, 0x13, 0x0B, 0x33, 0x2E, 0x1D, 0x13, 0x05, 0x1D,
	0x76, 0x54, 0x51, 0x2B, 0x0F, 0x03, 0x14, 0x37, 0x57, 0x2D, 0x0F, 0x5B,
	0x51, 0x21, 0x05, 0x1B, 0x01, 0x2F, 0x5C, 0x5C, 0x37, 0x1B, 0x28, 0x04,
	0x0A, 0x01, 0x16, 0x4E, 0x0C, 0x0A, 0x37, 0x5A, 0x25, 0x14, 0x3E, 0x08,
	0x59, 0x03, 0x18, 0x3C, 0x6D, 0x54, 0x32, 0x26, 0x1B, 0x13, 0x03, 0x07,
	0x29, 0x07, 0x20, 0x34, 0x20, 0x36, 0x0D, 0x0B, 0x36, 0x33, 0x5F, 0x3E,
	0x11, 0x59, 0x12, 0x26, 0x05, 0x26, 0x36, 0x58, 0x45, 0x44, 0x20, 0x3A,
	0x10, 0x05, 0x1D, 0x0A, 0x3C, 0x35, 0x07, 0x00, 0x26, 0x35, 0x32, 0x41,
	0x20, 0x3A, 0x5B, 0x2F, 0x1A, 0x24, 0x34, 0x3B, 0x57, 0x0B, 0x1F, 0x16,
	0x00, 0x16, 0x5A, 0x11, 0x09, 0x15, 0x06, 0x20, 0x07, 0x34, 0x1F, 0x30,
	0x1E, 0x5D, 0x2A, 0x09, 0x30, 0x14, 0x04, 0x27, 0x1E, 0x0E, 0x25, 0x5D,
	0x72, 0x1C, 0x29, 0x1E, 0x52, 0x0B, 0x5E, 0x0E, 0x3D, 0x5F, 0x21, 0x36,
	0x0E, 0x59, 0x5F, 0x32, 0x14, 0x08, 0x06, 0x0E, 0x26, 0x3E, 0x50, 0x03,
	0x01, 0x0E, 0x27, 0x10, 0x37, 0x5F, 0x3A, 0x05, 0x18, 0x1B, 0x33, 0x37,
	0x04, 0x2E, 0x1E, 0x5F, 0x15, 0x07, 0x18, 0x03, 0x5F, 0x69, 0x2A, 0x32,
	0x06, 0x1C, 0x75, 0x09, 0x02, 0x26, 0x1D, 0x0D, 0x47, 0x38, 0x36, 0x59,
	0x12, 0x2A, 0x2D, 0x3C, 0x05, 0x2D, 0x09, 0x0D, 0x17, 0x29, 0x18, 0x23,
	0x13, 0x0A, 0x5F, 0x0A, 0x54, 0x19, 0x1C, 0x44, 0x0D, 0x5F, 0x53, 0x19,
	0x5C, 0x00, 0x0A, 0x57, 0x37, 0x26, 0x17, 0x1A, 0x53, 0x2A, 0x13, 0x06,
	0x35, 0x39, 0x23, 0x26, 0x34, 0x07, 0x52, 0x22, 0x0E, 0x1A, 0x28, 0x54,
	0x5D, 0x5C, 0x23, 0x59, 0x0E, 0x1F, 0x5E, 0x77, 0x2D, 0x0D, 0x5E, 0x33,
	0x34, 0x1D, 0x56, 0x5A, 0x1B, 0x2F, 0x1A, 0x05, 0x59, 0x08, 0x27, 0x5F,
	0x13, 0x5B, 0x3D, 0x09, 0x24, 0x39, 0x0A, 0x33, 0x32, 0x2A, 0x10, 0x00,
	0x19, 0x70, 0x29, 0x05, 0x21, 0x05, 0x28, 0x28, 0x31, 0x1B, 0x3A, 0x12,
	0x3A, 0x2E, 0x5D, 0x2F, 0x12, 0x25, 0x34, 0x3E, 0x00, 0x7A, 0x3A, 0x11,
	0x0F, 0x0F, 0x38, 0x26, 0x09, 0x01, 0x03, 0x18, 0x54, 0x35, 0x0F, 0x1D,
	0x21, 0x09, 0x50, 0x04, 0x3D, 0x0A, 0x39, 0x4E, 0x1A, 0x12, 0x11, 0x1D,
	0x31, 0x3D, 0x05, 0x71, 0x0E, 0x4E, 0x02, 0x31, 0x6D, 0x1F, 0x32, 0x0A,
	0x3E, 0x04, 0x58, 0x14, 0x28, 0x5B, 0x0E, 0x5E, 0x4A, 0x17, 0x21, 0x0E,
	0x04, 0x4A, 0x03, 0x2F, 0x38, 0x34, 0x35, 0x05, 0x0D, 0x20, 0x2E, 0x3B,
	0x57, 0x33, 0x11, 0x35, 0x31, 0x1B, 0x02, 0x34, 0x5A, 0x28, 0x3E, 0x32,
	0x1A, 0x1D, 0x10, 0x0F, 0x23, 0x34, 0x36, 0x09, 0x57, 0x02, 0x6D, 0x58,
	0x12, 0x2B, 0x3F, 0x2A, 0x1B, 0x55, 0x14, 0x32, 0x32, 0x2F, 0x35, 0x56,
	0x13, 0x06, 0x16, 0x39, 0x04, 0x5C, 0x70, 0x0B, 0x08, 0x5B, 0x0E, 0x23,
	0x1D, 0x31, 0x0F, 0x03, 0x16, 0x2D, 0x07, 0x00, 0x3D, 0x24, 0x5D, 0x50,
	0x1A, 0x58, 0x6D, 0x22, 0x09, 0x5A, 0x13, 0x6D, 0x02, 0x23, 0x3A, 0x40,
	0x33, 0x0D, 0x26, 0x20, 0x26, 0x24, 0x5A, 0x2B, 0x45, 0x2A, 0x1A, 0x43,
	0x0D, 0x3E, 0x59, 0x01, 0x0A, 0x52, 0x34, 0x3D, 0x28, 0x3F, 0x52, 0x3D,
	0x03, 0x0C, 0x05, 0x0A, 0x38, 0x27, 0x18, 0x5B, 0x54, 0x29, 0x3E, 0x34,
	0x21, 0x4E, 0x05, 0x05, 0x6D, 0x0E, 0x35, 0x5C, 0x24, 0x17, 0x00, 0x05,
	0x34, 0x31, 0x24, 0x0E, 0x1B, 0x2C, 0x24, 0x32, 0x18, 0x17, 0x03, 0x00,
	0x35, 0x01, 0x03, 0x01, 0x08, 0x09, 0x25, 0x55, 0x3D, 0x3A, 0x26, 0x47,
	0x0D, 0x0A, 0x2C, 0x35, 0x05, 0x58, 0x0A, 0x28, 0x2E, 0x59, 0x03, 0x38,
	0x3E, 0x23, 0x09, 0x2C, 0x2D, 0x07, 0x0E, 0x03, 0x50, 0x28, 0x2F, 0x11,
	0x5A, 0x0B, 0x20, 0x3F, 0x3A, 0x3B, 0x4E, 0x1C, 0x44, 0x73, 0x25, 0x15,
	0x1B, 0x44, 0x3A, 0x2F, 0x2D, 0x0D, 0x0D, 0x69, 0x3D, 0x08, 0x5F, 0x27,
	0x24, 0x1F, 0x27, 0x04, 0x07, 0x74, 0x1C, 0x26, 0x2B, 0x1D, 0x38, 0x2B,
	0x0B, 0x2D, 0x03, 0x00, 0x02, 0x22, 0x3F, 0x39, 0x32, 0x5A, 0x39, 0x0C,
	0x5B, 0x28, 0x1E, 0x18, 0x45, 0x1C, 0x2F, 0x43, 0x34, 0x23, 0x1D, 0x6D,
	0x1E, 0x2E, 0x17, 0x5A, 0x2C, 0x5C, 0x27, 0x25, 0x0D, 0x7A, 0x24, 0x0C,
	0x1A, 0x1C, 0x33, 0x0E, 0x2B, 0x0B, 0x05, 0x2B, 0x06, 0x2F, 0x06, 0x3E,
	0x2F, 0x16, 0x30, 0x16, 0x1B, 0x71, 0x01, 0x26, 0x1A, 0x21, 0x20, 0x0E,
	0x1B, 0x25, 0x1D, 0x10, 0x24, 0x09, 0x09, 0x0E, 0x10, 0x09, 0x0F, 0x07,
	0x06, 0x12, 0x3E, 0x2A, 0x14, 0x1D, 0x71, 0x02, 0x26, 0x27, 0x01, 0x73,
	0x05, 0x02, 0x21, 0x00, 0x76, 0x1A, 0x0D, 0x37, 0x2E, 0x6D, 0x0D, 0x1B,
	0x3C, 0x03, 0x0D, 0x2E, 0x12, 0x39, 0x1D, 0x05, 0x36, 0x11, 0x0F, 0x5A,
	0x3A, 0x02, 0x04, 0x1B, 0x59, 0x17, 0x1B, 0x19, 0x23, 0x22, 0x07, 0x0F,
	0x3B, 0x06, 0x53, 0x35, 0x59, 0x35, 0x14, 0x59, 0x16, 0x27, 0x59, 0x0D,
	0x06, 0x05, 0x47, 0x02, 0x18, 0x24, 0x76, 0x2E, 0x55, 0x58, 0x21, 0x2B,
	0x14, 0x15, 0x04, 0x2A, 0x03, 0x19, 0x1B, 0x5B, 0x03, 0x27, 0x0A, 0x0F,
	0x1F, 0x40, 0x32, 0x1E, 0x22, 0x36, 0x5F, 0x05, 0x00, 0x14, 0x18, 0x2F,
	0x24, 0x5D, 0x23, 0x08, 0x07, 0x1A, 0x34, 0x2F, 0x29, 0x21, 0x2E, 0x3E,
	0x52, 0x3D, 0x3D, 0x07, 0x0E, 0x0A, 0x45, 0x44, 0x23, 0x05, 0x0F, 0x24,
	0x59, 0x75, 0x23, 0x31, 0x01, 0x01, 0x71, 0x5B, 0x37, 0x2B, 0x40, 0x0A,
	0x0D, 0x02, 0x56, 0x38, 0x10, 0x34, 0x17, 0x29, 0x24, 0x34, 0x3B, 0x13,
	0x58, 0x0F, 0x0A, 0x3C, 0x38, 0x5E, 0x0E, 0x33, 0x0E, 0x09, 0x18, 0x1A,
	0x2E, 0x2B, 0x2B, 0x3B, 0x19, 0x73, 0x1E, 0x59, 0x00, 0x3F, 0x14, 0x15,
	0x14, 0x0B, 0x22, 0x04, 0x5C, 0x0B, 0x58, 0x11, 0x12, 0x3E, 0x59, 0x2B,
	0x3F, 0x0E, 0x36, 0x3B, 0x5D, 0x0D, 0x0C, 0x59, 0x2C, 0x0B, 0x0C, 0x7A,
	0x22, 0x37, 0x23, 0x0E, 0x07, 0x5E, 0x32, 0x16, 0x18, 0x06, 0x5E, 0x54,
	0x3D, 0x3B, 0x1B, 0x39, 0x2E, 0x23, 0x1E, 0x27, 0x0A, 0x4A, 0x2C, 0x05,
	0x2A, 0x38, 0x50, 0x5F, 0x11, 0x07, 0x59, 0x1B, 0x28, 0x2F, 0x76, 0x5C,
	0x10, 0x0F, 0x5C, 0x06, 0x47, 0x29, 0x2D, 0x23, 0x73, 0x05, 0x59, 0x56,
	0x58, 0x3A, 0x27, 0x11, 0x5C, 0x04, 0x21, 0x2B, 0x37, 0x20, 0x33, 0x0B,
	0x3C, 0x51, 0x16, 0x0A, 0x7A, 0x59, 0x34, 0x0A, 0x11, 0x6D, 0x16, 0x07,
	0x29, 0x39, 0x0F, 0x21, 0x31, 0x58, 0x18, 0x27, 0x29, 0x51, 0x1E, 0x40,
	0x35, 0x3B, 0x38, 0x14, 0x03, 0x21, 0x5D, 0x55, 0x5C, 0x33, 0x36, 0x01,
	0x2C, 0x36, 0x0F, 0x15, 0x1A, 0x38, 0x45, 0x5B, 0x29, 0x22, 0x15, 0x0D,
	0x52, 0x7B, 0x01, 0x59, 0x1F, 0x07, 0x3B, 0x18, 0x32, 0x22, 0x1C, 0x15,
	0x1B, 0x39, 0x57, 0x0A, 0x0E, 0x18, 0x55, 0x18, 0x5A, 0x05, 0x01, 0x09,
	0x01, 0x00, 0x75, 0x5D, 0x10, 0x1B, 0x18, 0x35, 0x43, 0x32, 0x1A, 0x3B,
	0x7A, 0x0D, 0x16, 0x27, 0x0D, 0x2D, 0x08, 0x27, 0x17, 0x39, 0x74, 0x01,
	0x52, 0x1D, 0x1F, 0x69, 0x58, 0x37, 0x17, 0x2A, 0x2D, 0x00, 0x35, 0x59,
	0x5B, 0x08, 0x2A, 0x08, 0x36, 0x39, 0x73, 0x20, 0x24, 0x57, 0x0C, 0x71,
	0x25, 0x04, 0x06, 0x1F, 0x06, 0x1A, 0x0B, 0x3F, 0x03, 0x26, 0x22, 0x52,
	0x02, 0x0C, 0x0D, 0x38, 0x16, 0x29, 0x2C, 0x70, 0x2D, 0x22, 0x3E, 0x03,
	0x0F, 0x2D, 0x07, 0x19, 0x1A, 0x0C, 0x3B, 0x57, 0x59, 0x1D, 0x77, 0x5D,
	0x26, 0x5D, 0x39, 0x27, 0x18, 0x53, 0x0F, 0x3B, 0x29, 0x28, 0x4A, 0x2C,
	0x59, 0x15, 0x38, 0x23, 0x26, 0x00, 0x14, 0x22, 0x2D, 0x2C, 0x23, 0x33,
	0x0E, 0x00, 0x00, 0x08, 0x00, 0x5E, 0x34, 0x1E, 0x5F, 0x71, 0x26, 0x58,
	0x24, 0x59, 0x1A, 0x1A, 0x28, 0x22, 0x27, 0x09, 0x55, 0x30, 0x41, 0x1A,
	0x11, 0x5D, 0x24, 0x1B, 0x1C, 0x33, 0x01, 0x57, 0x2A, 0x07, 0x0C, 0x0A,
	0x36, 0x16, 0x3F, 0x73, 0x14, 0x00, 0x45, 0x1E, 0x35, 0x55, 0x35, 0x28,
	0x2F, 0x23, 0x5F, 0x00, 0x5D, 0x11, 0x71, 0x2E, 0x26, 0x5D, 0x5B, 0x1A,
	0x5A, 0x19, 0x08, 0x1A, 0x35, 0x1C, 0x37, 0x0A, 0x2D, 0x7A, 0x07, 0x19,
	0x59, 0x21, 0x36, 0x35, 0x37, 0x39, 0x3D, 0x34, 0x54, 0x51, 0x41, 0x5D,
	0x1B, 0x23, 0x53, 0x14, 0x19, 0x69, 0x16, 0x31, 0x18, 0x58, 0x03, 0x34,
	0x57, 0x16, 0x0F, 0x31, 0x55, 0x0D, 0x3E, 0x32, 0x28, 0x2A, 0x0D, 0x1C,
	0x38, 0x76, 0x5B, 0x2E, 0x3E, 0x5C, 0x01, 0x36, 0x4E, 0x19, 0x1D, 0x73,
	0x3A, 0x36, 0x38, 0x11, 0x36, 0x36, 0x59, 0x0A, 0x2D, 0x06, 0x36, 0x39,
	0x41, 0x04, 0x0E, 0x22, 0x2C, 0x3F, 0x1A, 0x20, 0x26, 0x35, 0x2A, 0x11,
	0x2B, 0x59, 0x24, 0x1F, 0x1D, 0x7B, 0x24, 0x13, 0x37, 0x02, 0x2F, 0x5F,
	0x14, 0x08, 0x09, 0x15, 0x27, 0x16, 0x3D, 0x0F, 0x17, 0x5E, 0x52, 0x37,
	0x19, 0x16, 0x0F, 0x00, 0x29, 0x27, 0x07, 0x3A, 0x0C, 0x56, 0x00, 0x07,
	0x1C, 0x0F, 0x5F, 0x09, 0x0C, 0x1C, 0x2C, 0x22, 0x11, 0x03, 0x0B, 0x2E,
	0x1D, 0x1C, 0x74, 0x35, 0x0A, 0x16, 0x11, 0x2F, 0x0E, 0x53, 0x2F, 0x12,
	0x70, 0x5B, 0x26, 0x34, 0x18, 0x7A, 0x2F, 0x12, 0x5B, 0x3F, 0x06, 0x3C,
	0x06, 0x39, 0x05, 0x15, 0x1A, 0x0D, 0x1F, 0x44, 0x17, 0x3C, 0x09, 0x5B,
	0x1D, 0x14, 0x1D, 0x50, 0x21, 0x13, 0x1A, 0x43, 0x16, 0x23, 0x53, 0x77,
	0x08, 0x03, 0x3F, 0x25, 0x27, 0x0E, 0x4A, 0x5A, 0x19, 0x69, 0x0B, 0x39,
	0x5F, 0x31, 0x27, 0x28, 0x0D, 0x41, 0x08, 0x0E, 0x3C, 0x36, 0x5F, 0x5E,
	0x34, 0x54, 0x20, 0x58, 0x1B, 0x36, 0x34, 0x51, 0x58, 0x2F, 0x36, 0x58,
	0x51, 0x0F, 0x19, 0x30, 0x27, 0x54, 0x21, 0x1A, 0x6D, 0x3A, 0x02, 0x29,
	0x1D, 0x0D, 0x01, 0x52, 0x05, 0x3C, 0x07, 0x55, 0x2E, 0x06, 0x5A, 0x7A,
	0x5F, 0x37, 0x59, 0x52, 0x12, 0x22, 0x08, 0x3B, 0x5B, 0x26, 0x2B, 0x0F,
	0x0A, 0x3C, 0x32, 0x47, 0x11, 0x1A, 0x38, 0x09, 0x5C, 0x35, 0x29, 0x0C,
	0x26, 0x0A, 0x20, 0x58, 0x1B, 0x29, 0x1C, 0x52, 0x00, 0x40, 0x16, 0x1A,
	0x17, 0x02, 0x05, 0x0E, 0x43, 0x37, 0x16, 0x52, 0x6D, 0x08, 0x50, 0x41,
	0x12, 0x7A, 0x55, 0x55, 0x0D, 0x59, 0x06, 0x1F, 0x2C, 0x0F, 0x21, 0x73,
	0x21, 0x0C, 0x18, 0x3E, 0x7A, 0x3B, 0x23, 0x5E, 0x5D, 0x0E, 0x21, 0x20,
	0x3E, 0x0D, 0x77, 0x39, 0x56, 0x16, 0x1F, 0x01, 0x3E, 0x12, 0x0B, 0x3A,
	0x73, 0x04, 0x0D, 0x08, 0x58, 0x10, 0x5B, 0x26, 0x14, 0x5A, 0x0F, 0x3A,
	0x07, 0x1F, 0x5C, 0x69, 0x1D, 0x13, 0x1B, 0x53, 0x75, 0x2F, 0x56, 0x39,
	0x44, 0x72, 0x59, 0x07, 0x1C, 0x02, 0x2D, 0x5B, 0x13, 0x56, 0x31, 0x3B,
	0x58, 0x35, 0x1C, 0x2D, 0x0C, 0x3F, 0x0C, 0x1C, 0x5B, 0x69, 0x35, 0x26,
	0x1A, 0x0F, 0x17, 0x1C, 0x13, 0x05, 0x07, 0x18, 0x02, 0x32, 0x58, 0x1E,
	0x0F, 0x3E, 0x52, 0x1D, 0x23, 0x6D, 0x01, 0x0E, 0x22, 0x26, 0x37, 0x1E,
	0x14, 0x02, 0x2C, 0x76, 0x5F, 0x0F, 0x28, 0x1F, 0x3B, 0x47, 0x0E, 0x0A,
	0x11, 0x72, 0x39, 0x50, 0x1F, 0x40, 0x2C, 0x0B, 0x14, 0x1D, 0x2A, 0x73,
	0x25, 0x2A, 0x1D, 0x27, 0x29, 0x14, 0x11, 0x1C, 0x01, 0x0E, 0x5A, 0x25,
	0x57, 0x1C, 0x34, 0x18, 0x04, 0x3D, 0x5C, 0x04, 0x1A, 0x07, 0x58, 0x38,
	0x38, 0x5D, 0x09, 0x1E, 0x05, 0x24, 0x43, 0x28, 0x14, 0x58, 0x1A, 0x0F,
	0x4A, 0x08, 0x40, 0x04, 0x0F, 0x03, 0x59, 0x02, 0x04, 0x5E, 0x1B, 0x21,
	0x3D, 0x7B, 0x05, 0x02, 0x22, 0x00, 0x70, 0x38, 0x11, 0x03, 0x32, 0x29,
	0x3E, 0x16, 0x5D, 0x01, 0x06, 0x26, 0x12, 0x2A, 0x59, 0x7A, 0x04, 0x15,
	0x1C, 0x05, 0x2C, 0x21, 0x0D, 0x23, 0x3D, 0x09, 0x3F, 0x0D, 0x22, 0x04,
	0x73, 0x2A, 0x23, 0x3D, 0x3B, 0x75, 0x20, 0x00, 0x3E, 0x38, 0x09, 0x01,
	0x11, 0x2D, 0x5D, 0x6D, 0x54, 0x0F, 0x18, 0x29, 0x0E, 0x58, 0x19, 0x0F,
	0x2A, 0x2E, 0x5F, 0x54, 0x1F, 0x2D, 0x14, 0x55, 0x23, 0x28, 0x28, 0x7A,
	0x3F, 0x00, 0x1F, 0x1F, 0x27, 0x01, 0x03, 0x28, 0x01, 0x73, 0x24, 0x15,
	0x1D, 0x3C, 0x72, 0x39, 0x04, 0x58, 0x5B, 0x05, 0x14, 0x3B, 0x0B, 0x05,
	0x74, 0x2A, 0x10, 0x39, 0x5C, 0x69, 0x38, 0x38, 0x1F, 0x1B, 0x74, 0x08,
	0x18, 0x00, 0x39, 0x35, 0x34, 0x10, 0x58, 0x04, 0x70, 0x1E, 0x52, 0x02,
	0x0A, 0x34, 0x5A, 0x11, 0x41, 0x3F, 0x27, 0x5B, 0x39, 0x41, 0x2D, 0x12,
	0x1E, 0x26, 0x5A, 0x0F, 0x31, 0x5D, 0x31, 0x5B, 0x27, 0x6D, 0x19, 0x4E,
	0x5A, 0x21, 0x6D, 0x1F, 0x39, 0x41, 0x2F, 0x12, 0x29, 0x00, 0x5B, 0x44,
	0x77, 0x23, 0x57, 0x06, 0x2C, 0x77, 0x34, 0x59, 0x25, 0x5A, 0x72, 0x3A,
	0x17, 0x45, 0x28, 0x24, 0x2F, 0x0E, 0x38, 0x44, 0x2A, 0x20, 0x39, 0x58,
	0x39, 0x6D, 0x2D, 0x17, 0x45, 0x3E, 0x24, 0x15, 0x22, 0x41, 0x5C, 0x08,
	0x47, 0x30, 0x36, 0x44, 0x2E, 0x3C, 0x53, 0x2D, 0x0D, 0x7A, 0x58, 0x13,
	0x41, 0x28, 0x0D, 0x05, 0x31, 0x5A, 0x0C, 0x2E, 0x38, 0x09, 0x00, 0x20,
	0x74, 0x34, 0x24, 0x24, 0x09, 0x14, 0x0B, 0x53, 0x5E, 0x5B, 0x35, 0x01,
	0x2C, 0x2A, 0x18, 0x17, 0x06, 0x2A, 0x24, 0x44, 0x70, 0x0D, 0x0A, 0x0B,
	0x38, 0x11, 0x25, 0x37, 0x41, 0x1B, 0x05, 0x43, 0x12, 0x5F, 0x59, 0x1A,
	0x0A, 0x57, 0x1C, 0x0D, 0x05, 0x36, 0x22, 0x36, 0x02, 0x6D, 0x0A, 0x4E,
	0x28, 0x3B, 0x21, 0x5E, 0x38, 0x28, 0x32, 0x26, 0x3A, 0x03, 0x1C, 0x1C,
	0x11, 0x39, 0x33, 0x28, 0x21, 0x1B, 0x1D, 0x2A, 0x07, 0x0C, 0x76, 0x5A,
	0x10, 0x25, 0x02, 0x2D, 0x2E, 0x31, 0x00, 0x1B, 0x29, 0x25, 0x54, 0x07,
	0x5E, 0x06, 0x09, 0x20, 0x2B, 0x04, 0x0E, 0x3D, 0x22, 0x3D, 0x38, 0x2B,
	0x01, 0x58, 0x3E, 0x05, 0x75, 0x23, 0x55, 0x45, 0x08, 0x12, 0x58, 0x55,
	0x0B, 0x5E, 0x7B, 0x19, 0x26, 0x1A, 0x2D, 0x2A, 0x29, 0x15, 0x3D, 0x04,
	0x05, 0x2A, 0x27, 0x3C, 0x2E, 0x76, 0x22, 0x2A, 0x2A, 0x20, 0x0F, 0x14,
	0x30, 0x3D, 0x33, 0x09, 0x14, 0x28, 0x16, 0x02, 0x25, 0x05, 0x2E, 0x04,
	0x2C, 0x11, 0x43, 0x0B, 0x5A, 0x22, 0x25, 0x23, 0x2A, 0x05, 0x31, 0x05,
	0x2B, 0x04, 0x3B, 0x5D, 0x28, 0x21, 0x00, 0x27, 0x33, 0x36, 0x3F, 0x0E,
	0x5D, 0x5A, 0x30, 0x5D, 0x12, 0x5D, 0x0E, 0x36, 0x09, 0x17, 0x08, 0x1B,
	0x08, 0x1A, 0x14, 0x59, 0x11, 0x73, 0x15, 0x04, 0x3C, 0x52, 0x12, 0x55,
	0x58, 0x1F, 0x19, 0x7B, 0x5B, 0x11, 0x45, 0x1A, 0x14, 0x3B, 0x14, 0x1A,
	0x3C, 0x30, 0x3B, 0x10, 0x3E, 0x3B, 0x32, 0x16, 0x52, 0x08, 0x3A, 0x76,
	0x55, 0x56, 0x18, 0x11, 0x0C, 0x07, 0x06, 0x45, 0x31, 0x33, 0x5D, 0x3B,
	0x1A, 0x23, 0x0E, 0x1A, 0x04, 0x27, 0x06, 0x7B, 0x59, 0x59, 0x59, 0x3C,
	0x73, 0x1B, 0x05, 0x24, 0x5E, 0x32, 0x2F, 0x37, 0x25, 0x3A, 0x11, 0x22,
	0x14, 0x07, 0x04, 0x7B, 0x21, 0x26, 0x45, 0x2C, 0x23, 0x15, 0x31, 0x1A,
	0x21, 0x18, 0x01, 0x00, 0x3F, 0x2F, 0x77, 0x3C, 0x18, 0x2B, 0x24, 0x28,
	0x14, 0x27, 0x18, 0x40, 0x2C, 0x3B, 0x35, 0x5C, 0x02, 0x04, 0x35, 0x4E,
	0x27, 0x0E, 0x11, 0x35, 0x30, 0x26, 0x5E, 0x0E, 0x15, 0x25, 0x0C, 0x5C,
	0x3A, 0x04, 0x35, 0x17, 0x59, 0x09, 0x07, 0x57, 0x05, 0x11, 0x36, 0x2A,
	0x0F, 0x05, 0x23, 0x0B, 0x38, 0x0E, 0x29, 0x53, 0x2B, 0x26, 0x20, 0x57,
	0x2A, 0x32, 0x00, 0x25, 0x17, 0x25, 0x76, 0x29, 0x12, 0x0F, 0x0E, 0x0E,
	0x43, 0x37, 0x06, 0x1C, 0x0E, 0x09, 0x27, 0x39, 0x22, 0x7B, 0x15, 0x1B,
	0x0F, 0x3D, 0x10, 0x58, 0x52, 0x05, 0x12, 0x71, 0x3A, 0x38, 0x02, 0x0A,
	0x38, 0x36, 0x0E, 0x24, 0x06, 0x28, 0x0E, 0x11, 0x2D, 0x32, 0x36, 0x26,
	0x56, 0x2A, 0x05, 0x3B, 0x5A, 0x54, 0x07, 0x0E, 0x72, 0x29, 0x19, 0x58,
	0x1C, 0x30, 0x0D, 0x22, 0x00, 0x05, 0x72, 0x08, 0x26, 0x0C, 0x1E, 0x33,
	0x09, 0x23, 0x5A, 0x01, 0x18, 0x3B, 0x12, 0x17, 0x3E, 0x25, 0x36, 0x30,
	0x16, 0x04, 0x3B, 0x39, 0x52, 0x3D, 0x3B, 0x1B, 0x04, 0x58, 0x37, 0x33,
	0x12, 0x1C, 0x13, 0x5A, 0x1C, 0x2A, 0x0B, 0x07, 0x5A, 0x05, 0x7A, 0x1D,
	0x54, 0x04, 0x07, 0x11, 0x1E, 0x56, 0x20, 0x0A, 0x26, 0x27, 0x00, 0x08,
	0x22, 0x6D, 0x3E, 0x30, 0x56, 0x1E, 0x20, 0x04, 0x14, 0x34, 0x22, 0x7A,
	0x07, 0x27, 0x23, 0x3F, 0x6D, 0x3E, 0x18, 0x37, 0x3E, 0x70, 0x3C, 0x58,
	0x26, 0x20, 0x04, 0x14, 0x0B, 0x41, 0x2D, 0x38, 0x04, 0x2F, 0x59, 0x5B,
	0x0C, 0x28, 0x4A, 0x5D, 0x5E, 0x69, 0x36, 0x02, 0x59, 0x20, 0x27, 0x2E,
	0x4E, 0x3F, 0x12, 0x35, 0x38, 0x16, 0x2A, 0x59, 0x13, 0x3B, 0x25, 0x08,
	0x00, 0x76, 0x1A, 0x58, 0x2A, 0x27, 0x01, 0x0A, 0x23, 0x08, 0x31, 0x08,
	0x1B, 0x29, 0x5A, 0x01, 0x31, 0x22, 0x4A, 0x3C, 0x02, 0x6D, 0x5C, 0x09,
	0x37, 0x23, 0x7A, 0x29, 0x53, 0x25, 0x08, 0x03, 0x47, 0x55, 0x0B, 0x2A,
	0x24, 0x34, 0x59, 0x1B, 0x52, 0x30, 0x3C, 0x20, 0x3E, 0x1E, 0x1B, 0x26,
	0x31, 0x18, 0x18, 0x72, 0x35, 0x31, 0x56, 0x18, 0x31, 0x22, 0x4A, 0x0C,
	0x02, 0x6D, 0x5C, 0x02, 0x1D, 0x22, 0x7A, 0x28, 0x58, 0x07, 0x5E, 0x25,
	0x3C, 0x16, 0x04, 0x18, 0x2A, 0x5F, 0x2A, 0x16, 0x3B, 0x35, 0x20, 0x12,
	0x2B, 0x5F, 0x00, 0x55, 0x2D, 0x1C, 0x29, 0x6D, 0x29, 0x58, 0x09, 0x0D,
	0x3B, 0x21, 0x37, 0x0B, 0x0E, 0x0E, 0x0E, 0x31, 0x3E, 0x0C, 0x2C, 0x35,
	0x27, 0x19, 0x23, 0x75, 0x0F, 0x36, 0x2F, 0x44, 0x2F, 0x03, 0x15, 0x57,
	0x2F, 0x0E, 0x2E, 0x31, 0x2F, 0x0D, 0x20, 0x00, 0x16, 0x26, 0x5F, 0x23,
	0x5E, 0x28, 0x41, 0x05, 0x1B, 0x04, 0x59, 0x22, 0x5C, 0x0C, 0x23, 0x20,
	0x18, 0x3A, 0x24, 0x35, 0x1B, 0x19, 0x23, 0x75, 0x15, 0x37, 0x14, 0x18,
	0x76, 0x58, 0x22, 0x57, 0x28, 0x7B, 0x06, 0x39, 0x2F, 0x0D, 0x34, 0x06,
	0x0F, 0x1B, 0x5D, 0x38, 0x02, 0x59, 0x59, 0x2D, 0x12, 0x04, 0x56, 0x37,
	0x5E, 0x35, 0x26, 0x56, 0x29, 0x0F, 0x25, 0x02, 0x20, 0x3E, 0x1F, 0x06,
	0x19, 0x05, 0x09, 0x05, 0x03, 0x3C, 0x12, 0x07, 0x32, 0x09, 0x54, 0x22,
	0x45, 0x13, 0x10, 0x0B, 0x31, 0x5B, 0x0E, 0x0E, 0x0A, 0x32, 0x25, 0x1C,
	0x0E, 0x1B, 0x07, 0x5C, 0x2C, 0x0C, 0x05, 0x56, 0x09, 0x09, 0x72, 0x1B,
	0x2A, 0x19, 0x44, 0x75, 0x26, 0x26, 0x2A, 0x1D, 0x03, 0x0A, 0x00, 0x1A,
	0x1C, 0x0E, 0x58, 0x2A, 0x5C, 0x26, 0x24, 0x01, 0x38, 0x1E, 0x53, 0x01,
	0x5B, 0x26, 0x38, 0x0C, 0x71, 0x58, 0x26, 0x14, 0x2F, 0x0E, 0x2F, 0x31,
	0x14, 0x53, 0x17, 0x47, 0x27, 0x0A, 0x02, 0x30, 0x1B, 0x2D, 0x5A, 0x27,
	0x18, 0x14, 0x0D, 0x09, 0x05, 0x77, 0x05, 0x2D, 0x08, 0x39, 0x33, 0x1B,
	0x19, 0x56, 0x28, 0x69, 0x2B, 0x58, 0x09, 0x44, 0x03, 0x09, 0x18, 0x3A,
	0x08, 0x75, 0x24, 0x31, 0x2F, 0x3B, 0x23, 0x18, 0x16, 0x22, 0x5F, 0x1A,
	0x5E, 0x20, 0x56, 0x2A, 0x69, 0x55, 0x33, 0x0D, 0x5C, 0x04, 0x5F, 0x20,
	0x18, 0x03, 0x71, 0x35, 0x58, 0x19, 0x23, 0x75, 0x0A, 0x02, 0x2F, 0x40,
	0x0B, 0x14, 0x05, 0x59, 0x25, 0x75, 0x28, 0x17, 0x2F, 0x3B, 0x1B, 0x28,
	0x16, 0x3E, 0x5F, 0x03, 0x1F, 0x29, 0x08, 0x05, 0x1B, 0x1C, 0x59, 0x22,
	0x5C, 0x0E, 0x19, 0x20, 0x41, 0x38, 0x01, 0x1B, 0x29, 0x19, 0x3B, 0x70,
	0x09, 0x03, 0x00, 0x32, 0x77, 0x1B, 0x29, 0x59, 0x09, 0x2F, 0x2D, 0x4E,
	0x2A, 0x24, 0x35, 0x3C, 0x20, 0x18, 0x1D, 0x11, 0x34, 0x2E, 0x17, 0x27,
	0x25, 0x24, 0x51, 0x18, 0x18, 0x00, 0x43, 0x23, 0x21, 0x3A, 0x75, 0x35,
	0x37, 0x45, 0x31, 0x2B, 0x34, 0x16, 0x1C, 0x18, 0x69, 0x58, 0x25, 0x57,
	0x2C, 0x0E, 0x2E, 0x1B, 0x16, 0x38, 0x16, 0x26, 0x17, 0x04, 0x32, 0x1A,
	0x47, 0x52, 0x24, 0x0C, 0x12, 0x1B, 0x25, 0x1D, 0x21, 0x76, 0x28, 0x58,
	0x16, 0x08, 0x01, 0x47, 0x31, 0x06, 0x0D, 0x75, 0x3F, 0x0C, 0x2F, 0x44,
	0x01, 0x23, 0x18, 0x00, 0x0C, 0x0E, 0x5C, 0x2D, 0x5C, 0x2A, 0x26, 0x15,
	0x12, 0x08, 0x08, 0x03, 0x47, 0x53, 0x28, 0x0C, 0x12, 0x1B, 0x31, 0x1D,
	0x02, 0x76, 0x2F, 0x58, 0x03, 0x32, 0x36, 0x55, 0x2D, 0x0C, 0x2A, 0x24,
	0x2D, 0x07, 0x0F, 0x11, 0x35, 0x20, 0x55, 0x2D, 0x59, 0x06, 0x0A, 0x0F,
	0x37, 0x07, 0x7A, 0x24, 0x56, 0x23, 0x0E, 0x03, 0x43, 0x33, 0x28, 0x0C,
	0x1A, 0x1B, 0x17, 0x1D, 0x59, 0x71, 0x27, 0x19, 0x1C, 0x1C, 0x24, 0x5E,
	0x24, 0x56, 0x2A, 0x69, 0x36, 0x0E, 0x14, 0x3B, 0x71, 0x0B, 0x17, 0x1D,
	0x25, 0x69, 0x36, 0x08, 0x22, 0x1C, 0x12, 0x5B, 0x2A, 0x39, 0x2A, 0x24,
	0x2E, 0x4A, 0x16, 0x3D, 0x1B, 0x22, 0x4A, 0x34, 0x02, 0x71, 0x5C, 0x20,
	0x5C, 0x26, 0x7A, 0x2D, 0x4A, 0x19, 0x39, 0x25, 0x24, 0x16, 0x3A, 0x59,
	0x2F, 0x5F, 0x2E, 0x16, 0x3D, 0x76, 0x24, 0x58, 0x22, 0x27, 0x00, 0x3C,
	0x20, 0x18, 0x09, 0x30, 0x0B, 0x39, 0x5F, 0x3B, 0x0E, 0x1A, 0x38, 0x03,
	0x18, 0x06, 0x54, 0x22, 0x59, 0x2D, 0x0D, 0x2D, 0x07, 0x3C, 0x0E, 0x35,
	0x5F, 0x54, 0x29, 0x27, 0x12, 0x3D, 0x03, 0x5C, 0x26, 0x17, 0x54, 0x24,
	0x2A, 0x13, 0x30, 0x35, 0x31, 0x19, 0x09, 0x31, 0x47, 0x52, 0x21, 0x13,
	0x20, 0x1B, 0x03, 0x5C, 0x08, 0x21, 0x28, 0x04, 0x2C, 0x0E, 0x3A, 0x5F,
	0x20, 0x18, 0x1E, 0x7B, 0x19, 0x05, 0x07, 0x58, 0x03, 0x1A, 0x12, 0x2B,
	0x32, 0x08, 0x54, 0x2D, 0x59, 0x2E, 0x27, 0x2D, 0x4E, 0x38, 0x2A, 0x37,
	0x55, 0x0C, 0x5D, 0x04, 0x13, 0x3D, 0x31, 0x59, 0x22, 0x2F, 0x2D, 0x4E,
	0x2F, 0x40, 0x35, 0x3C, 0x54, 0x29, 0x27, 0x24, 0x06, 0x09, 0x5A, 0x5B,
	0x31, 0x2F, 0x59, 0x26, 0x52, 0x2C, 0x3C, 0x20, 0x08, 0x01, 0x13, 0x34,
	0x4A, 0x5A, 0x58, 0x2D, 0x3D, 0x30, 0x20, 0x5C, 0x06, 0x5B, 0x23, 0x14,
	0x09, 0x10, 0x1E, 0x31, 0x08, 0x53, 0x6D, 0x2A, 0x17, 0x09, 0x26, 0x7B,
	0x0D, 0x26, 0x2C, 0x0D, 0x00, 0x47, 0x16, 0x3A, 0x0C, 0x12, 0x5D, 0x0A,
	0x22, 0x1D, 0x23, 0x08, 0x57, 0x2B, 0x2E, 0x06, 0x09, 0x19, 0x00, 0x32,
	0x08, 0x1B, 0x29, 0x59, 0x5D, 0x14, 0x16, 0x12, 0x1B, 0x52, 0x01, 0x28,
	0x23, 0x18, 0x32, 0x33, 0x1F, 0x2D, 0x56, 0x32, 0x70, 0x2E, 0x4E, 0x25,
	0x13, 0x1A, 0x58, 0x1B, 0x0B, 0x1F, 0x06, 0x2D, 0x29, 0x09, 0x3B, 0x75,
	0x08, 0x26, 0x2F, 0x44, 0x2E, 0x58, 0x15, 0x57, 0x25, 0x71, 0x1E, 0x30,
	0x19, 0x27, 0x76, 0x3A, 0x53, 0x2D, 0x53, 0x0A, 0x55, 0x12, 0x22, 0x18,
	0x12, 0x23, 0x19, 0x59, 0x0C, 0x0A, 0x5C, 0x05, 0x1D, 0x2C, 0x7A, 0x24,
	0x58, 0x18, 0x33, 0x03, 0x3C, 0x0B, 0x37, 0x33, 0x69, 0x5D, 0x56, 0x5E,
	0x58, 0x76, 0x2A, 0x58, 0x2C, 0x5C, 0x03, 0x5F, 0x06, 0x36, 0x5A, 0x7A,
	0x20, 0x17, 0x37, 0x5C, 0x72, 0x24, 0x59, 0x26, 0x52, 0x2E, 0x5F, 0x20,
	0x18, 0x0C, 0x1A, 0x35, 0x2B, 0x45, 0x31, 0x2B, 0x5F, 0x55, 0x08, 0x40,
	0x0D, 0x5B, 0x25, 0x18, 0x29, 0x34, 0x0E, 0x15, 0x41, 0x5E, 0x24, 0x35,
	0x58, 0x58, 0x3B, 0x6D, 0x28, 0x14, 0x16, 0x5C, 0x25, 0x0A, 0x51, 0x03,
	0x32, 0x08, 0x47, 0x02, 0x07, 0x44, 0x72, 0x2D, 0x4A, 0x1B, 0x44, 0x03,
	0x1A, 0x06, 0x41, 0x32, 0x12, 0x1B, 0x2D, 0x1D, 0x3E, 0x71, 0x23, 0x19,
	0x5D, 0x5F, 0x34, 0x47, 0x2E, 0x59, 0x2A, 0x24, 0x2D, 0x31, 0x34, 0x3B,
	0x03, 0x1A, 0x14, 0x23, 0x33, 0x0D, 0x1B, 0x29, 0x5E, 0x33, 0x7A, 0x24,
	0x58, 0x01, 0x3B, 0x03, 0x1A, 0x09, 0x41, 0x32, 0x37, 0x5F, 0x2E, 0x16,
	0x23, 0x72, 0x20, 0x4E, 0x26, 0x0F, 0x25, 0x3C, 0x20, 0x41, 0x1E, 0x1A,
	0x0B, 0x29, 0x5F, 0x0E, 0x0E, 0x1A, 0x03, 0x2A, 0x5D, 0x0E, 0x54, 0x25,
	0x45, 0x13, 0x04, 0x0B, 0x4E, 0x14, 0x1A, 0x35, 0x20, 0x59, 0x5D, 0x2D,
	0x6D, 0x0B, 0x25, 0x58, 0x5C, 0x7A, 0x2E, 0x4A, 0x2A, 0x25, 0x28, 0x43,
	0x25, 0x0A, 0x03, 0x1A, 0x59, 0x0C, 0x27, 0x44, 0x25, 0x1A, 0x55, 0x59,
	0x18, 0x08, 0x54, 0x20, 0x57, 0x0C, 0x27, 0x2E, 0x07, 0x39, 0x5B, 0x37,
	0x55, 0x10, 0x3E, 0x04, 0x34, 0x1B, 0x31, 0x59, 0x20, 0x15, 0x28, 0x4E,
	0x2C, 0x09, 0x01, 0x1A, 0x1B, 0x56, 0x3D, 0x69, 0x28, 0x31, 0x5F, 0x58,
	0x1B, 0x28, 0x59, 0x2A, 0x5C, 0x0E, 0x54, 0x25, 0x57, 0x04, 0x04, 0x0F,
	0x56, 0x23, 0x0D, 0x10, 0x0A, 0x16, 0x08, 0x59, 0x31, 0x54, 0x23, 0x0B,
	0x0E, 0x09, 0x0E, 0x31, 0x5D, 0x18, 0x38, 0x2A, 0x07, 0x09, 0x27, 0x7B,
	0x08, 0x53, 0x2C, 0x44, 0x00, 0x22, 0x0B, 0x26, 0x2A, 0x24, 0x1A, 0x0C,
	0x36, 0x24, 0x35, 0x02, 0x51, 0x36, 0x53, 0x0A, 0x08, 0x10, 0x59, 0x3F,
	0x08, 0x08, 0x0A, 0x00, 0x2A, 0x34, 0x19, 0x53, 0x36, 0x24, 0x3B, 0x02,
	0x51, 0x26, 0x53, 0x0A, 0x55, 0x0F, 0x26, 0x2A, 0x12, 0x04, 0x0F, 0x37,
	0x09, 0x7A, 0x16, 0x27, 0x08, 0x03, 0x30, 0x55, 0x05, 0x5C, 0x28, 0x24,
	0x2D, 0x2E, 0x16, 0x3F, 0x25, 0x34, 0x50, 0x00, 0x27, 0x34, 0x35, 0x1B,
	0x58, 0x27, 0x7A, 0x28, 0x4A, 0x17, 0x39, 0x25, 0x02, 0x16, 0x26, 0x18,
	0x0C, 0x47, 0x05, 0x07, 0x0D, 0x35, 0x06, 0x58, 0x0A, 0x59, 0x01, 0x0A,
	0x20, 0x1B, 0x12, 0x34, 0x2E, 0x31, 0x37, 0x52, 0x37, 0x08, 0x0B, 0x3E,
	0x04, 0x34, 0x43, 0x4A, 0x24, 0x21, 0x7B, 0x55, 0x26, 0x1C, 0x2A, 0x34,
	0x2D, 0x31, 0x37, 0x5C, 0x21, 0x1E, 0x26, 0x08, 0x3A, 0x6D, 0x54, 0x05,
	0x5C, 0x27, 0x37, 0x2D, 0x07, 0x3A, 0x06, 0x35, 0x5B, 0x59, 0x41, 0x2D,
	0x6D, 0x0B, 0x0B, 0x58, 0x5C, 0x7A, 0x2D, 0x4A, 0x28, 0x52, 0x2A, 0x5B,
	0x06, 0x3E, 0x58, 0x27, 0x34, 0x2E, 0x17, 0x08, 0x2F, 0x23, 0x31, 0x5B,
	0x5C, 0x7A, 0x2F, 0x4A, 0x2D, 0x25, 0x28, 0x0A, 0x23, 0x21, 0x12, 0x0A,
	0x0F, 0x13, 0x29, 0x3B, 0x03, 0x0A, 0x38, 0x1E, 0x1C, 0x0E, 0x58, 0x02,
	0x5C, 0x2A, 0x27, 0x2D, 0x4E, 0x37, 0x2D, 0x21, 0x5B, 0x26, 0x21, 0x29,
	0x24, 0x3E, 0x10, 0x19, 0x52, 0x35, 0x2E, 0x56, 0x2B, 0x52, 0x2B, 0x3C,
	0x54, 0x03, 0x22, 0x24, 0x2E, 0x4A, 0x16, 0x0F, 0x35, 0x20, 0x55, 0x21,
	0x59, 0x06, 0x0F, 0x25, 0x45, 0x44, 0x04, 0x0F, 0x56, 0x21, 0x24, 0x00,
	0x0A, 0x32, 0x58, 0x1C, 0x2E, 0x58, 0x27, 0x57, 0x2C, 0x75, 0x2F, 0x07,
	0x14, 0x26, 0x17, 0x47, 0x20, 0x0A, 0x0C, 0x1A, 0x2D, 0x39, 0x1D, 0x3D,
	0x70, 0x22, 0x59, 0x28, 0x5C, 0x09, 0x08, 0x1B, 0x1D, 0x3E, 0x7A, 0x29,
	0x58, 0x1B, 0x33, 0x03, 0x24, 0x06, 0x3E, 0x5C, 0x69, 0x58, 0x29, 0x57,
	0x04, 0x14, 0x16, 0x12, 0x05, 0x5F, 0x01, 0x55, 0x23, 0x57, 0x02, 0x71,
	0x2D, 0x17, 0x1A, 0x23, 0x25, 0x3C, 0x50, 0x0D, 0x27, 0x34, 0x0E, 0x2B,
	0x19, 0x27, 0x76, 0x23, 0x53, 0x22, 0x08, 0x06, 0x47, 0x50, 0x5B, 0x0C,
	0x0E, 0x5F, 0x35, 0x02, 0x3C, 0x2C, 0x54, 0x29, 0x57, 0x01, 0x09, 0x1B,
	0x56, 0x19, 0x2F, 0x70, 0x0A, 0x02, 0x2F, 0x40, 0x0C, 0x04, 0x07, 0x59,
	0x3D, 0x05, 0x2F, 0x17, 0x2F, 0x1D, 0x31, 0x19, 0x38, 0x22, 0x53, 0x0A,
	0x5E, 0x2C, 0x08, 0x05, 0x1B, 0x1C, 0x59, 0x29, 0x5C, 0x06, 0x2B, 0x16,
	0x59, 0x1C, 0x20, 0x5E, 0x30, 0x56, 0x2A, 0x69, 0x21, 0x33, 0x08, 0x5C,
	0x06, 0x2B, 0x25, 0x08, 0x28, 0x37, 0x14, 0x56, 0x09, 0x0D, 0x70, 0x0E,
	0x16, 0x2A, 0x5F, 0x77, 0x2A, 0x52, 0x1D, 0x33, 0x31, 0x2B, 0x59, 0x26,
	0x52, 0x2C, 0x5F, 0x20, 0x08, 0x0C, 0x38, 0x35, 0x11, 0x45, 0x31, 0x2B,
	0x02, 0x16, 0x18, 0x18, 0x37, 0x58, 0x25, 0x57, 0x22, 0x0E, 0x2F, 0x07,
	0x2C, 0x1D, 0x1B, 0x36, 0x14, 0x0A, 0x0C, 0x1A, 0x2D, 0x07, 0x1A, 0x0E,
	0x1B, 0x28, 0x59, 0x2D, 0x5C, 0x0B, 0x54, 0x20, 0x0B, 0x58, 0x21, 0x19,
	0x58, 0x1F, 0x33, 0x03, 0x1A, 0x06, 0x41, 0x32, 0x28, 0x1B, 0x29, 0x59,
	0x5F, 0x77, 0x5B, 0x0D, 0x1D, 0x53, 0x6D, 0x20, 0x19, 0x0C, 0x5F, 0x11,
	0x5E, 0x20, 0x56, 0x28, 0x69, 0x15, 0x0F, 0x5E, 0x21, 0x2D, 0x2E, 0x58,
	0x0F, 0x38, 0x75, 0x5E, 0x29, 0x03, 0x2A, 0x6D, 0x28, 0x2E, 0x16, 0x05,
	0x25, 0x3C, 0x51, 0x28, 0x1C, 0x0E, 0x58, 0x18, 0x28, 0x44, 0x36, 0x0D,
	0x38, 0x2A, 0x53, 0x01, 0x5B, 0x26, 0x0B, 0x29, 0x24, 0x3E, 0x10, 0x19,
	0x19, 0x7A, 0x5F, 0x27, 0x18, 0x0C, 0x75, 0x35, 0x0B, 0x19, 0x23, 0x75,
	0x25, 0x59, 0x2F, 0x40, 0x00, 0x55, 0x0B, 0x36, 0x5E, 0x70, 0x26, 0x07,
	0x2A, 0x40, 0x35, 0x02, 0x06, 0x26, 0x59, 0x0F, 0x34, 0x4E, 0x57, 0x1C,
	0x38, 0x06, 0x19, 0x09, 0x23, 0x7A, 0x06, 0x27, 0x36, 0x0C, 0x20, 0x5E,
	0x34, 0x56, 0x2A, 0x69, 0x28, 0x15, 0x07, 0x33, 0x03, 0x5F, 0x12, 0x14,
	0x2D, 0x6D, 0x1F, 0x20, 0x1D, 0x21, 0x7A, 0x2E, 0x58, 0x09, 0x05, 0x03,
	0x0A, 0x06, 0x5C, 0x1C, 0x20, 0x54, 0x56, 0x28, 0x33, 0x25, 0x34, 0x53,
	0x1D, 0x53, 0x03, 0x47, 0x22, 0x0A, 0x01, 0x1A, 0x1C, 0x4A, 0x16, 0x06,
	0x71, 0x54, 0x35, 0x1B, 0x13, 0x76, 0x5D, 0x04, 0x34, 0x11, 0x0E, 0x22,
	0x33, 0x0C, 0x0F, 0x73, 0x26, 0x11, 0x5F, 0x53, 0x26, 0x3E, 0x12, 0x26,
	0x18, 0x07, 0x55, 0x19, 0x3F, 0x3A, 0x0A, 0x47, 0x16, 0x36, 0x25, 0x2E,
	0x15, 0x3B, 0x14, 0x3B, 0x0E, 0x0B, 0x25, 0x57, 0x2D, 0x0E, 0x23, 0x0C,
	0x28, 0x0C, 0x38, 0x5B, 0x22, 0x26, 0x3E, 0x2F, 0x25, 0x39, 0x41, 0x0E,
	0x38, 0x0E, 0x24, 0x5D, 0x11, 0x71, 0x5B, 0x0F, 0x2D, 0x26, 0x6D, 0x47,
	0x4E, 0x45, 0x28, 0x77, 0x19, 0x10, 0x0F, 0x26, 0x1A, 0x07, 0x31, 0x17,
	0x00, 0x29, 0x09, 0x04, 0x20, 0x20, 0x30, 0x21, 0x11, 0x3B, 0x58, 0x20,
	0x22, 0x51, 0x0F, 0x04, 0x0F, 0x54, 0x0F, 0x34, 0x5A, 0x69, 0x58, 0x4A,
	0x1D, 0x18, 0x28, 0x08, 0x33, 0x5C, 0x31, 0x69, 0x5C, 0x02, 0x56, 0x40,
	0x7A, 0x06, 0x57, 0x1E, 0x52, 0x12, 0x5E, 0x59, 0x1C, 0x1F, 0x00, 0x1C,
	0x0F, 0x5F, 0x3F, 0x74, 0x0A, 0x12, 0x0F, 0x02, 0x38, 0x27, 0x31, 0x37,
	0x44, 0x1A, 0x24, 0x10, 0x3E, 0x3B, 0x18, 0x26, 0x0B, 0x36, 0x58, 0x2B,
	0x5A, 0x31, 0x1B, 0x00, 0x06, 0x1C, 0x52, 0x26, 0x11, 0x2D, 0x5A, 0x0B,
	0x23, 0x28, 0x2D, 0x59, 0x09, 0x5D, 0x13, 0x17, 0x1D, 0x19, 0x1A, 0x33,
	0x38, 0x3F, 0x20, 0x59, 0x32, 0x28, 0x1A, 0x0A, 0x5B, 0x25, 0x13, 0x04,
	0x25, 0x45, 0x5A, 0x76, 0x20, 0x17, 0x34, 0x1E, 0x72, 0x2D, 0x0A, 0x59,
	0x3A, 0x01, 0x0F, 0x02, 0x09, 0x27, 0x2C, 0x0B, 0x30, 0x08, 0x3F, 0x73,
	0x0F, 0x13, 0x26, 0x3B, 0x03, 0x43, 0x03, 0x0A, 0x1C, 0x0A, 0x58, 0x38,
	0x5C, 0x29, 0x7B, 0x2B, 0x39, 0x17, 0x53, 0x1A, 0x47, 0x52, 0x24, 0x0C,
	0x12, 0x1B, 0x25, 0x1D, 0x21, 0x76, 0x28, 0x58, 0x17, 0x0A, 0x01, 0x22,
	0x29, 0x56, 0x19, 0x04, 0x0A, 0x09, 0x3C, 0x59, 0x0C, 0x14, 0x16, 0x0C,
	0x5D, 0x75, 0x21, 0x4E, 0x0D, 0x1A, 0x0A, 0x3C, 0x17, 0x09, 0x1B, 0x3B,
	0x5B, 0x2C, 0x41, 0x07, 0x1B, 0x06, 0x59, 0x2D, 0x5C, 0x07, 0x09, 0x20,
	0x41, 0x38, 0x3B, 0x1B, 0x1B, 0x19, 0x33, 0x70, 0x1B, 0x08, 0x38, 0x5E,
	0x70, 0x2E, 0x59, 0x2F, 0x52, 0x31, 0x3C, 0x20, 0x08, 0x0C, 0x20, 0x35,
	0x39, 0x19, 0x11, 0x31, 0x35, 0x52, 0x21, 0x13, 0x0A, 0x1B, 0x03, 0x5C,
	0x0C, 0x7A, 0x2E, 0x4A, 0x2D, 0x1F, 0x2B, 0x0A, 0x22, 0x0B, 0x11, 0x28,
	0x0F, 0x56, 0x2B, 0x0D, 0x03, 0x1A, 0x38, 0x2A, 0x1C, 0x0A, 0x58, 0x22,
	0x5C, 0x26, 0x21, 0x2D, 0x4A, 0x56, 0x39, 0x21, 0x5B, 0x20, 0x0B, 0x29,
	0x24, 0x3E, 0x4A, 0x19, 0x23, 0x35, 0x3C, 0x53, 0x5D, 0x11, 0x72, 0x3A,
	0x07, 0x22, 0x5A, 0x21, 0x5B, 0x31, 0x0D, 0x28, 0x69, 0x5D, 0x54, 0x09,
	0x3B, 0x35, 0x20, 0x12, 0x3E, 0x1C, 0x12, 0x5E, 0x10, 0x0C, 0x05, 0x1B,
	0x28, 0x16, 0x2A, 0x5C, 0x20, 0x01, 0x20, 0x41, 0x2F, 0x0D, 0x16, 0x29,
	0x09, 0x33, 0x73, 0x2B, 0x2D, 0x18, 0x09, 0x7B, 0x1B, 0x2D, 0x5A, 0x27,
	0x70, 0x2D, 0x59, 0x2D, 0x40, 0x70, 0x2A, 0x06, 0x59, 0x53, 0x75, 0x2A,
	0x17, 0x09, 0x44, 0x1B, 0x08, 0x16, 0x2A, 0x5C, 0x03, 0x3B, 0x25, 0x41,
	0x29, 0x0E, 0x28, 0x31, 0x17, 0x53, 0x14, 0x47, 0x23, 0x59, 0x29, 0x34,
	0x2E, 0x4E, 0x34, 0x52, 0x35, 0x3C, 0x54, 0x45, 0x32, 0x04, 0x47, 0x00,
	0x07, 0x58, 0x72, 0x1A, 0x12, 0x29, 0x53, 0x04, 0x55, 0x13, 0x5D, 0x2A,
	0x6D, 0x05, 0x54, 0x09, 0x33, 0x77, 0x01, 0x2D, 0x08, 0x3A, 0x69, 0x1B,
	0x19, 0x56, 0x28, 0x69, 0x2B, 0x58, 0x07, 0x19, 0x35, 0x20, 0x55, 0x5C,
	0x2D, 0x6D, 0x18, 0x14, 0x37, 0x20, 0x7A, 0x2F, 0x4A, 0x17, 0x5E, 0x25,
	0x34, 0x16, 0x08, 0x18, 0x74, 0x5F, 0x2E, 0x16, 0x58, 0x35, 0x16, 0x12,
	0x34, 0x3C, 0x06, 0x0A, 0x20, 0x0B, 0x12, 0x0E, 0x0B, 0x29, 0x5E, 0x0C,
	0x04, 0x43, 0x12, 0x1B, 0x32, 0x04, 0x54, 0x29, 0x59, 0x25, 0x37, 0x2E,
	0x07, 0x3C, 0x0A, 0x35, 0x22, 0x52, 0x21, 0x13, 0x75, 0x1B, 0x35, 0x5C,
	0x23, 0x2F, 0x28, 0x07, 0x2D, 0x1E, 0x3B, 0x38, 0x06, 0x26, 0x5A, 0x38,
	0x20, 0x17, 0x37, 0x0F, 0x35, 0x20, 0x55, 0x0D, 0x59, 0x05, 0x22, 0x06,
	0x08, 0x12, 0x09, 0x1B, 0x03, 0x56, 0x1D, 0x04, 0x0A, 0x08, 0x21, 0x1C,
	0x0E, 0x1B, 0x2D, 0x5C, 0x20, 0x30, 0x28, 0x4E, 0x37, 0x09, 0x38, 0x3C,
	0x07, 0x03, 0x26, 0x37, 0x55, 0x14, 0x5D, 0x2A, 0x12, 0x04, 0x07, 0x37,
	0x12, 0x38, 0x06, 0x2D, 0x2F, 0x3B, 0x34, 0x23, 0x39, 0x21, 0x11, 0x20,
	0x0B, 0x2D, 0x5E, 0x27, 0x70, 0x22, 0x02, 0x2C, 0x40, 0x35, 0x47, 0x20,
	0x41, 0x0E, 0x18, 0x0F, 0x56, 0x28, 0x1E, 0x00, 0x0A, 0x33, 0x1F, 0x1C,
	0x7B, 0x1B, 0x25, 0x59, 0x25, 0x76, 0x2A, 0x58, 0x3A, 0x12, 0x75, 0x5E,
	0x1B, 0x0D, 0x2A, 0x69, 0x2E, 0x05, 0x07, 0x33, 0x03, 0x43, 0x15, 0x00,
	0x0C, 0x24, 0x5E, 0x2E, 0x36, 0x24, 0x35, 0x14, 0x12, 0x2B, 0x53, 0x01,
	0x55, 0x0A, 0x36, 0x2A, 0x34, 0x0B, 0x17, 0x37, 0x52, 0x69, 0x08, 0x08,
	0x0C, 0x40, 0x08, 0x19, 0x3B, 0x39, 0x28, 0x24, 0x2F, 0x4A, 0x14, 0x09,
	0x25, 0x0A, 0x52, 0x0B, 0x33, 0x0D, 0x14, 0x37, 0x5D, 0x20, 0x29, 0x22,
	0x56, 0x28, 0x58, 0x03, 0x34, 0x06, 0x08, 0x59, 0x13, 0x5B, 0x0F, 0x37,
	0x29, 0x71, 0x2F, 0x39, 0x21, 0x19, 0x00, 0x3C, 0x20, 0x41, 0x32, 0x71,
	0x2D, 0x07, 0x1D, 0x2F, 0x37, 0x08, 0x0B, 0x22, 0x1E, 0x07, 0x3C, 0x4E,
	0x56, 0x3F, 0x75, 0x5B, 0x27, 0x29, 0x29, 0x24, 0x2D, 0x04, 0x16, 0x23,
	0x21, 0x5B, 0x26, 0x18, 0x13, 0x69, 0x03, 0x24, 0x19, 0x2F, 0x76, 0x26,
	0x53, 0x21, 0x08, 0x03, 0x47, 0x4E, 0x28, 0x08, 0x75, 0x23, 0x14, 0x2F,
	0x44, 0x13, 0x15, 0x16, 0x3A, 0x1C, 0x06, 0x5E, 0x27, 0x19, 0x2F, 0x75,
	0x15, 0x37, 0x14, 0x18, 0x23, 0x58, 0x29, 0x57, 0x2D, 0x0E, 0x2F, 0x31,
	0x2F, 0x44, 0x20, 0x24, 0x20, 0x08, 0x1D, 0x32, 0x34, 0x2E, 0x19, 0x52,
	0x35, 0x24, 0x55, 0x2D, 0x59, 0x0F, 0x0F, 0x20, 0x45, 0x5C, 0x2F, 0x02,
	0x4A, 0x21, 0x1C, 0x12, 0x59, 0x36, 0x24, 0x0D, 0x2B, 0x0A, 0x55, 0x59,
	0x18, 0x06, 0x55, 0x18, 0x09, 0x08, 0x6D, 0x47, 0x22, 0x5C, 0x2A, 0x6D,
	0x00, 0x55, 0x1A, 0x52, 0x0D, 0x0A, 0x13, 0x18, 0x1C, 0x0A, 0x58, 0x36,
	0x5C, 0x23, 0x7A, 0x2D, 0x56, 0x26, 0x13, 0x25, 0x15, 0x00, 0x20, 0x05,
	0x1A, 0x58, 0x13, 0x45, 0x24, 0x75, 0x2F, 0x07, 0x2F, 0x0D, 0x23, 0x1A,
	0x20, 0x41, 0x1D, 0x1B, 0x34, 0x2E, 0x17, 0x27, 0x72, 0x24, 0x59, 0x26,
	0x52, 0x2E, 0x3C, 0x20, 0x18, 0x0C, 0x6D, 0x35, 0x19, 0x45, 0x0F, 0x2B,
	0x02, 0x55, 0x08, 0x40, 0x0D, 0x5B, 0x22, 0x08, 0x2A, 0x12, 0x0E, 0x05,
	0x19, 0x2F, 0x76, 0x14, 0x27, 0x41, 0x1F, 0x21, 0x55, 0x2F, 0x45, 0x29,
	0x6D, 0x3E, 0x08, 0x19, 0x5C, 0x35, 0x28, 0x53, 0x17, 0x09, 0x2C, 0x35,
	0x14, 0x57, 0x2D, 0x6D, 0x2E, 0x4E, 0x37, 0x01, 0x35, 0x20, 0x55, 0x28,
	0x59, 0x09, 0x0A, 0x0C, 0x37, 0x1E, 0x7B, 0x2F, 0x4E, 0x16, 0x58, 0x1B,
	0x28, 0x16, 0x3E, 0x5C, 0x03, 0x20, 0x25, 0x3E, 0x12, 0x0F, 0x39, 0x4A,
	0x2F, 0x44, 0x73, 0x5F, 0x38, 0x2A, 0x53, 0x0B, 0x5B, 0x25, 0x5D, 0x2A,
	0x71, 0x1C, 0x53, 0x22, 0x0D, 0x10, 0x1E, 0x57, 0x59, 0x53, 0x00, 0x47,
	0x20, 0x20, 0x0C, 0x34, 0x2E, 0x4E, 0x34, 0x5E, 0x37, 0x08, 0x08, 0x00,
	0x04, 0x34, 0x54, 0x2E, 0x59, 0x3B, 0x37, 0x2D, 0x07, 0x3D, 0x1A, 0x35,
	0x20, 0x59, 0x5D, 0x2D, 0x12, 0x0B, 0x39, 0x57, 0x0F, 0x70, 0x28, 0x07,
	0x2D, 0x40, 0x35, 0x38, 0x06, 0x36, 0x5A, 0x2E, 0x20, 0x17, 0x0C, 0x21,
	0x74, 0x20, 0x59, 0x2A, 0x40, 0x70, 0x59, 0x06, 0x26, 0x1C, 0x12, 0x1F,
	0x00, 0x5D, 0x24, 0x3A, 0x38, 0x51, 0x22, 0x44, 0x0A, 0x08, 0x09, 0x5D,
	0x2A, 0x24, 0x1A, 0x11, 0x24, 0x44, 0x34, 0x1F, 0x57, 0x5D, 0x24, 0x3A,
	0x38, 0x51, 0x3A, 0x44, 0x0A, 0x08, 0x09, 0x5D, 0x2A, 0x12, 0x19, 0x4E,
	0x2F, 0x0D, 0x36, 0x2D, 0x2D, 0x18, 0x32, 0x08, 0x5A, 0x2D, 0x56, 0x2F,
	0x69, 0x5F, 0x3B, 0x09, 0x1D, 0x35, 0x43, 0x38, 0x03, 0x5C, 0x2C, 0x35,
	0x19, 0x58, 0x3B, 0x6D, 0x28, 0x14, 0x16, 0x09, 0x25, 0x0A, 0x51, 0x21,
	0x32, 0x0C, 0x47, 0x02, 0x07, 0x58, 0x72, 0x0F, 0x4A, 0x1B, 0x44, 0x03,
	0x24, 0x06, 0x3E, 0x5C, 0x16, 0x0F, 0x22, 0x45, 0x27, 0x10, 0x0A, 0x56,
	0x39, 0x3B, 0x16, 0x0A, 0x06, 0x0C, 0x5B, 0x09, 0x5B, 0x25, 0x29, 0x1C,
	0x71, 0x59, 0x08, 0x22, 0x0D, 0x13, 0x16, 0x57, 0x59, 0x53, 0x00, 0x09,
	0x23, 0x18, 0x32, 0x71, 0x2D, 0x07, 0x18, 0x24, 0x1A, 0x23, 0x16, 0x28,
	0x52, 0x0C, 0x47, 0x23, 0x08, 0x39, 0x70, 0x1B, 0x17, 0x16, 0x09, 0x1B,
	0x0E, 0x59, 0x59, 0x2D, 0x6D, 0x0B, 0x08, 0x0D, 0x29, 0x16, 0x07, 0x2F,
	0x5C, 0x23, 0x37, 0x2D, 0x07, 0x3F, 0x5D, 0x35, 0x5B, 0x59, 0x00, 0x2D,
	0x24, 0x0B, 0x56, 0x37, 0x1B, 0x35, 0x28, 0x56, 0x0D, 0x06, 0x01, 0x0A,
	0x25, 0x21, 0x13, 0x71, 0x59, 0x26, 0x27, 0x44, 0x01, 0x47, 0x18, 0x3A,
	0x0C, 0x0A, 0x5C, 0x33, 0x1D, 0x2F, 0x7A, 0x36, 0x53, 0x3E, 0x0D, 0x2C,
	0x35, 0x0F, 0x56, 0x22, 0x70, 0x2F, 0x02, 0x2F, 0x40, 0x73, 0x14, 0x06,
	0x41, 0x53, 0x0C, 0x2A, 0x31, 0x18, 0x1E, 0x7B, 0x19, 0x05, 0x04, 0x3B,
	0x03, 0x3C, 0x12, 0x5A, 0x32, 0x0D, 0x54, 0x22, 0x57, 0x0C, 0x27, 0x2E,
	0x4E, 0x38, 0x2A, 0x37, 0x55, 0x15, 0x3E, 0x2A, 0x12, 0x0B, 0x03, 0x37,
	0x1B, 0x35, 0x24, 0x56, 0x3B, 0x3C, 0x00, 0x43, 0x28, 0x2C, 0x0D, 0x75,
	0x27, 0x36, 0x2C, 0x44, 0x00, 0x21, 0x55, 0x41, 0x05, 0x13, 0x20, 0x12,
	0x57, 0x1C, 0x06, 0x5B, 0x51, 0x38, 0x11, 0x31, 0x26, 0x55, 0x26, 0x52,
	0x0E, 0x20, 0x23, 0x3E, 0x2A, 0x34, 0x0D, 0x58, 0x19, 0x23, 0x76, 0x54,
	0x27, 0x41, 0x18, 0x08, 0x35, 0x25, 0x56, 0x2F, 0x75, 0x2E, 0x2E, 0x2F,
	0x0D, 0x10, 0x09, 0x16, 0x00, 0x53, 0x38, 0x2A, 0x07, 0x06, 0x11, 0x1B,
	0x38, 0x16, 0x26, 0x5C, 0x0D, 0x2B, 0x22, 0x41, 0x23, 0x36, 0x04, 0x31,
	0x5B, 0x59, 0x0B, 0x43, 0x23, 0x1B, 0x1C, 0x2C, 0x0B, 0x29, 0x5E, 0x26,
	0x31, 0x2D, 0x59, 0x2D, 0x40, 0x72, 0x23, 0x54, 0x5C, 0x22, 0x7A, 0x2F,
	0x4A, 0x14, 0x2D, 0x25, 0x0A, 0x57, 0x3F, 0x2A, 0x31, 0x1B, 0x18, 0x19,
	0x05, 0x7A, 0x1A, 0x27, 0x08, 0x0C, 0x16, 0x35, 0x0B, 0x19, 0x2F, 0x75,
	0x3B, 0x36, 0x2C, 0x0D, 0x03, 0x23, 0x18, 0x28, 0x38, 0x71, 0x23, 0x15,
	0x18, 0x1C, 0x12, 0x5B, 0x38, 0x39, 0x2A, 0x6D, 0x2D, 0x4A, 0x16, 0x0F,
	0x35, 0x28, 0x55, 0x5C, 0x2D, 0x6D, 0x18, 0x09, 0x37, 0x2F, 0x7A, 0x25,
	0x56, 0x25, 0x0E, 0x03, 0x0A, 0x33, 0x25, 0x1C, 0x28, 0x54, 0x4E, 0x28,
	0x0D, 0x25, 0x06, 0x38, 0x2A, 0x1C, 0x06, 0x5B, 0x22, 0x39, 0x29, 0x6D,
	0x25, 0x13, 0x2C, 0x3B, 0x38, 0x21, 0x37, 0x45, 0x2E, 0x0C, 0x06, 0x52,
	0x2F, 0x0D, 0x31, 0x14, 0x38, 0x26, 0x52, 0x76, 0x02, 0x2C, 0x56, 0x40,
	0x0D, 0x3E, 0x07, 0x59, 0x1D, 0x21, 0x2F, 0x4A, 0x28, 0x52, 0x2B, 0x3C,
	0x20, 0x3E, 0x18, 0x32, 0x35, 0x2B, 0x45, 0x0A, 0x2B, 0x43, 0x51, 0x2F,
	0x18, 0x0D, 0x54, 0x26, 0x57, 0x18, 0x12, 0x2D, 0x07, 0x09, 0x11, 0x1B,
	0x36, 0x4A, 0x3C, 0x02, 0x71, 0x1B, 0x4E, 0x1D, 0x1E, 0x76, 0x28, 0x58,
	0x27, 0x27, 0x06, 0x0A, 0x23, 0x45, 0x11, 0x26, 0x19, 0x05, 0x04, 0x58,
	0x03, 0x0A, 0x12, 0x21, 0x32, 0x06, 0x54, 0x20, 0x59, 0x3B, 0x37, 0x2D,
	0x07, 0x38, 0x5F, 0x37, 0x55, 0x0B, 0x1B, 0x2A, 0x24, 0x38, 0x14, 0x19,
	0x5C, 0x35, 0x3C, 0x53, 0x04, 0x1C, 0x0A, 0x5B, 0x51, 0x02, 0x11, 0x31,
	0x09, 0x55, 0x28, 0x52, 0x09, 0x5B, 0x25, 0x18, 0x29, 0x24, 0x35, 0x05,
	0x19, 0x27, 0x76, 0x15, 0x27, 0x41, 0x18, 0x27, 0x35, 0x28, 0x45, 0x29,
	0x24, 0x38, 0x04, 0x19, 0x1D, 0x3A, 0x34, 0x38, 0x5F, 0x40, 0x18, 0x05,
	0x52, 0x19, 0x58, 0x31, 0x3A, 0x36, 0x2A, 0x0D, 0x00, 0x09, 0x19, 0x20,
	0x32, 0x04, 0x47, 0x07, 0x07, 0x44, 0x73, 0x01, 0x38, 0x2D, 0x53, 0x06,
	0x47, 0x16, 0x5B, 0x0C, 0x1A, 0x1B, 0x07, 0x1D, 0x2A, 0x75, 0x02, 0x38,
	0x0A, 0x1C, 0x0A, 0x5B, 0x2E, 0x03, 0x2F, 0x24, 0x28, 0x14, 0x19, 0x19,
	0x25, 0x0E, 0x53, 0x34, 0x02, 0x71, 0x5C, 0x0F, 0x1D, 0x3B, 0x21, 0x2D,
	0x4A, 0x5F, 0x31, 0x25, 0x34, 0x16, 0x2A, 0x18, 0x2F, 0x5F, 0x2E, 0x16,
	0x5C, 0x35, 0x28, 0x53, 0x5B, 0x08, 0x03, 0x09, 0x20, 0x41, 0x1E, 0x17,
	0x00, 0x2F, 0x5D, 0x00, 0x71, 0x20, 0x56, 0x09, 0x28, 0x23, 0x3C, 0x0F,
	0x39, 0x1A, 0x24, 0x34, 0x12, 0x0C, 0x05, 0x15, 0x28, 0x11, 0x0B, 0x25,
	0x03, 0x55, 0x08, 0x00, 0x1E, 0x09, 0x2D, 0x20, 0x41, 0x40, 0x01, 0x59,
	0x12, 0x03, 0x3A, 0x27, 0x3E, 0x00, 0x59, 0x5A, 0x00, 0x24, 0x12, 0x41,
	0x22, 0x69, 0x3E, 0x00, 0x19, 0x5C, 0x0D, 0x5B, 0x56, 0x56, 0x0E, 0x27,
	0x2F, 0x25, 0x0C, 0x28, 0x31, 0x43, 0x59, 0x41, 0x0E, 0x09, 0x5A, 0x14,
	0x23, 0x3F, 0x1B, 0x20, 0x05, 0x5A, 0x39, 0x21, 0x0D, 0x1B, 0x58, 0x29,
	0x23, 0x14, 0x32, 0x34, 0x38, 0x76, 0x43, 0x3B, 0x2D, 0x2E, 0x0C, 0x3B,
	0x13, 0x1C, 0x33, 0x6D, 0x34, 0x28, 0x56, 0x1E, 0x7B, 0x1B, 0x20, 0x17,
	0x3C, 0x31, 0x09, 0x2C, 0x56, 0x58, 0x34, 0x08, 0x2F, 0x23, 0x01, 0x35,
	0x5F, 0x16, 0x2F, 0x31, 0x6D, 0x03, 0x17, 0x3E, 0x04, 0x7B, 0x09, 0x0D,
	0x5F, 0x5C, 0x05, 0x55, 0x03, 0x09, 0x12, 0x0F, 0x02, 0x3B, 0x5D, 0x44,
	0x25, 0x5B, 0x50, 0x1B, 0x09, 0x2F, 0x24, 0x51, 0x36, 0x0C, 0x24, 0x3C,
	0x56, 0x1C, 0x5F, 0x24, 0x54, 0x4A, 0x17, 0x19, 0x38, 0x5A, 0x31, 0x36,
	0x44, 0x13, 0x54, 0x4A, 0x38, 0x5A, 0x24, 0x34, 0x04, 0x39, 0x3F, 0x76,
	0x06, 0x19, 0x1D, 0x58, 0x27, 0x1D, 0x4E, 0x0C, 0x05, 0x2F, 0x38, 0x55,
	0x34, 0x5E, 0x35, 0x39, 0x03, 0x24, 0x5E, 0x7B, 0x3D, 0x4E, 0x22, 0x18,
	0x32, 0x09, 0x27, 0x45, 0x3B, 0x2A, 0x20, 0x0E, 0x5A, 0x07, 0x0B, 0x1E,
	0x25, 0x1B, 0x1F, 0x2E, 0x27, 0x56, 0x0A, 0x1B, 0x33, 0x1A, 0x55, 0x18,
	0x05, 0x6D, 0x27, 0x0B, 0x5D, 0x44, 0x06, 0x0A, 0x24, 0x22, 0x27, 0x6D,
	0x39, 0x11, 0x5D, 0x11, 0x2C, 0x43, 0x0A, 0x3B, 0x44, 0x76, 0x22, 0x17,
	0x04, 0x3B, 0x7A, 0x18, 0x26, 0x21, 0x3B, 0x21, 0x35, 0x38, 0x0A, 0x3F,
	0x0A, 0x38, 0x4A, 0x3F, 0x58, 0x06, 0x3C, 0x2D, 0x0D, 0x24, 0x1B, 0x43,
	0x39, 0x1B, 0x1C, 0x70, 0x07, 0x0F, 0x05, 0x04, 0x70, 0x38, 0x14, 0x3F,
	0x0D, 0x18, 0x5F, 0x58, 0x24, 0x2F, 0x0C, 0x04, 0x0D, 0x22, 0x5B, 0x06,
	0x55, 0x54, 0x3E, 0x26, 0x03, 0x1B, 0x0F, 0x36, 0x59, 0x07, 0x1B, 0x14,
	0x0A, 0x09, 0x32, 0x03, 0x10, 0x28, 0x1F, 0x2C, 0x5B, 0x32, 0x41, 0x0C,
	0x24, 0x5C, 0x07, 0x23, 0x06, 0x6D, 0x43, 0x2D, 0x36, 0x44, 0x13, 0x5B,
	0x2A, 0x06, 0x39, 0x69, 0x38, 0x06, 0x06, 0x23, 0x2F, 0x43, 0x0D, 0x1A,
	0x33, 0x04, 0x0B, 0x28, 0x09, 0x18, 0x70, 0x00, 0x38, 0x27, 0x18, 0x69,
	0x3B, 0x04, 0x1D, 0x21, 0x00, 0x3F, 0x17, 0x14, 0x1E, 0x74, 0x0A, 0x56,
	0x1C, 0x31, 0x75, 0x58, 0x34, 0x06, 0x52, 0x77, 0x3C, 0x08, 0x2F, 0x11,
	0x03, 0x3A, 0x0D, 0x2F, 0x02, 0x06, 0x5F, 0x50, 0x3F, 0x28, 0x0C, 0x1A,
	0x23, 0x24, 0x00, 0x00, 0x3D, 0x2D, 0x37, 0x2F, 0x7A, 0x01, 0x27, 0x2D,
	0x21, 0x32, 0x18, 0x13, 0x0F, 0x24, 0x10, 0x47, 0x0A, 0x3E, 0x00, 0x15,
	0x25, 0x25, 0x56, 0x2E, 0x77, 0x2B, 0x04, 0x2F, 0x44, 0x03, 0x2B, 0x30,
	0x28, 0x5C, 0x75, 0x21, 0x33, 0x5F, 0x5C, 0x73, 0x1F, 0x0B, 0x3C, 0x3C,
	0x2D, 0x26, 0x26, 0x38, 0x22, 0x04, 0x21, 0x24, 0x34, 0x29, 0x0F, 0x0B,
	0x2F, 0x19, 0x18, 0x29, 0x5A, 0x20, 0x41, 0x01, 0x18, 0x1D, 0x36, 0x0D,
	0x5A, 0x0F, 0x0E, 0x34, 0x23, 0x05, 0x27, 0x38, 0x1B, 0x2D, 0x27, 0x3A,
	0x14, 0x06, 0x59, 0x2F, 0x26, 0x34, 0x55, 0x2B, 0x12, 0x0F, 0x54, 0x2B,
	0x1D, 0x0D, 0x15, 0x06, 0x2F, 0x3E, 0x21, 0x20, 0x3D, 0x15, 0x0F, 0x09,
	0x34, 0x1D, 0x26, 0x3C, 0x28, 0x11, 0x54, 0x17, 0x28, 0x24, 0x3B, 0x0D,
	0x13, 0x5E, 0x31, 0x27, 0x54, 0x0F, 0x24, 0x5C, 0x31, 0x1F, 0x3B, 0x05,
	0x0C, 0x7A, 0x14, 0x57, 0x1B, 0x33, 0x6D, 0x00, 0x18, 0x19, 0x2C, 0x77,
	0x2A, 0x11, 0x2D, 0x29, 0x2E, 0x5A, 0x04, 0x16, 0x3E, 0x76, 0x5C, 0x2C,
	0x09, 0x53, 0x35, 0x22, 0x0B, 0x25, 0x13, 0x73, 0x5B, 0x4A, 0x08, 0x3F,
	0x0B, 0x3C, 0x2C, 0x3E, 0x0C, 0x00, 0x1B, 0x23, 0x5B, 0x20, 0x27, 0x2D,
	0x4E, 0x2F, 0x5D, 0x13, 0x14, 0x51, 0x5D, 0x11, 0x29, 0x0D, 0x02, 0x2A,
	0x26, 0x2A, 0x5E, 0x30, 0x45, 0x32, 0x01, 0x54, 0x0F, 0x1E, 0x2D, 0x18,
	0x5B, 0x17, 0x18, 0x31, 0x13, 0x21, 0x08, 0x5C, 0x0A, 0x7B, 0x5E, 0x0F,
	0x5C, 0x2A, 0x15, 0x18, 0x56, 0x07, 0x39, 0x29, 0x16, 0x4A, 0x56, 0x1E,
	0x0C, 0x23, 0x2E, 0x22, 0x44, 0x71, 0x5C, 0x05, 0x34, 0x2E, 0x76, 0x2D,
	0x59, 0x07, 0x1F, 0x03, 0x0A, 0x0A, 0x41, 0x22, 0x01, 0x0A, 0x27, 0x20,
	0x23, 0x71, 0x19, 0x19, 0x22, 0x44, 0x0C, 0x54, 0x30, 0x21, 0x32, 0x0B,
	0x26, 0x26, 0x5B, 0x2E, 0x1A, 0x35, 0x36, 0x2D, 0x27, 0x71, 0x21, 0x37,
	0x17, 0x3D, 0x2A, 0x0E, 0x30, 0x07, 0x26, 0x20, 0x58, 0x35, 0x1C, 0x1D,
	0x00, 0x23, 0x35, 0x04, 0x0C, 0x0C, 0x1B, 0x27, 0x17, 0x25, 0x21, 0x25,
	0x36, 0x34, 0x0D, 0x72, 0x5F, 0x0A, 0x1E, 0x58, 0x0F, 0x2E, 0x23, 0x1B,
	0x52, 0x2F, 0x3B, 0x2E, 0x05, 0x5F, 0x35, 0x55, 0x0A, 0x5E, 0x22, 0x28,
	0x43, 0x16, 0x36, 0x33, 0x69, 0x36, 0x2F, 0x2C, 0x52, 0x0A, 0x04, 0x39,
	0x21, 0x53, 0x16, 0x0B, 0x2A, 0x0D, 0x31, 0x0C, 0x1C, 0x53, 0x1A, 0x0F,
	0x74, 0x1A, 0x00, 0x58, 0x1D, 0x3B, 0x25, 0x0A, 0x28, 0x01, 0x73, 0x54,
	0x27, 0x07, 0x23, 0x75, 0x26, 0x56, 0x1E, 0x5D, 0x1B, 0x43, 0x54, 0x5E,
	0x44, 0x38, 0x1D, 0x13, 0x2F, 0x0A, 0x29, 0x2D, 0x59, 0x00, 0x31, 0x03,
	0x5F, 0x06, 0x08, 0x22, 0x1A, 0x35, 0x25, 0x0D, 0x28, 0x7A, 0x04, 0x52,
	0x2D, 0x27, 0x05, 0x09, 0x0D, 0x2B, 0x31, 0x69, 0x2D, 0x35, 0x25, 0x2D,
	0x14, 0x43, 0x0B, 0x27, 0x39, 0x1B, 0x28, 0x2C, 0x2C, 0x06, 0x13, 0x09,
	0x28, 0x21, 0x53, 0x03, 0x24, 0x39, 0x5A, 0x07, 0x3B, 0x26, 0x30, 0x2F,
	0x59, 0x13, 0x0E, 0x28, 0x14, 0x32, 0x06, 0x0F, 0x32, 0x0D, 0x03, 0x74,
	0x5C, 0x02, 0x23, 0x3B, 0x01, 0x59, 0x0D, 0x29, 0x2D, 0x03, 0x3E, 0x25,
	0x16, 0x0E, 0x32, 0x2B, 0x53, 0x0B, 0x1B, 0x24, 0x3F, 0x36, 0x0C, 0x2C,
	0x26, 0x09, 0x56, 0x37, 0x24, 0x13, 0x08, 0x39, 0x08, 0x1D, 0x3B, 0x21,
	0x2F, 0x2D, 0x5E, 0x74, 0x35, 0x00, 0x28, 0x1D, 0x16, 0x00, 0x02, 0x3F,
	0x13, 0x23, 0x5D, 0x4A, 0x25, 0x0D, 0x12, 0x54, 0x26, 0x36, 0x5D, 0x30,
	0x3A, 0x16, 0x20, 0x12, 0x0C, 0x3F, 0x20, 0x06, 0x22, 0x05, 0x47, 0x03,
	0x05, 0x3C, 0x20, 0x01, 0x00, 0x45, 0x3A, 0x70, 0x07, 0x31, 0x05, 0x26,
	0x0B, 0x2D, 0x02, 0x2C, 0x40, 0x11, 0x35, 0x06, 0x16, 0x1C, 0x06, 0x59,
	0x56, 0x37, 0x13, 0x72, 0x06, 0x02, 0x20, 0x53, 0x72, 0x59, 0x0C, 0x45,
	0x11, 0x05, 0x14, 0x20, 0x02, 0x0C, 0x0F, 0x3F, 0x20, 0x18, 0x22, 0x15,
	0x3D, 0x29, 0x37, 0x29, 0x7A, 0x00, 0x0D, 0x2F, 0x23, 0x2B, 0x28, 0x24,
	0x38, 0x0C, 0x13, 0x15, 0x2C, 0x45, 0x1C, 0x0E, 0x0A, 0x3B, 0x00, 0x1D,
	0x13, 0x1D, 0x14, 0x3A, 0x0C, 0x05, 0x15, 0x57, 0x17, 0x2E, 0x26, 0x47,
	0x25, 0x14, 0x27, 0x12, 0x01, 0x04, 0x3B, 0x01, 0x31, 0x1B, 0x08, 0x34,
	0x27, 0x0A, 0x1E, 0x22, 0x29, 0x5B, 0x01, 0x01, 0x32, 0x0D, 0x0C, 0x2A,
	0x21, 0x37, 0x45, 0x53, 0x0A, 0x5E, 0x35, 0x1B, 0x2A, 0x37, 0x3D, 0x13,
	0x09, 0x3B, 0x35, 0x16, 0x28, 0x2A, 0x53, 0x04, 0x59, 0x27, 0x0B, 0x2E,
	0x2C, 0x2E, 0x26, 0x0F, 0x52, 0x25, 0x54, 0x06, 0x0D, 0x52, 0x04, 0x1F,
	0x29, 0x5B, 0x00, 0x0B, 0x15, 0x24, 0x1D, 0x2A, 0x27, 0x3D, 0x51, 0x06,
	0x3B, 0x17, 0x25, 0x0B, 0x1C, 0x38, 0x1A, 0x07, 0x0A, 0x3B, 0x3F, 0x75,
	0x39, 0x04, 0x56, 0x24, 0x15, 0x5A, 0x50, 0x29, 0x12, 0x69, 0x5A, 0x28,
	0x5F, 0x11, 0x08, 0x55, 0x02, 0x24, 0x5B, 0x26, 0x0B, 0x29, 0x19, 0x2E,
	0x29, 0x29, 0x59, 0x2A, 0x53, 0x28, 0x3A, 0x22, 0x5A, 0x00, 0x16, 0x0E,
	0x51, 0x28, 0x13, 0x13, 0x1F, 0x31, 0x45, 0x08, 0x30, 0x5C, 0x16, 0x17,
	0x31, 0x7A, 0x3B, 0x1B, 0x41, 0x1C, 0x11, 0x19, 0x02, 0x19, 0x5D, 0x13,
	0x1F, 0x37, 0x5E, 0x40, 0x7A, 0x00, 0x19, 0x2D, 0x12, 0x31, 0x26, 0x14,
	0x58, 0x38, 0x18, 0x07, 0x0C, 0x1A, 0x2F, 0x38, 0x15, 0x57, 0x2A, 0x3D,
	0x73, 0x35, 0x25, 0x5E, 0x2E, 0x38, 0x26, 0x26, 0x1A, 0x25, 0x2D, 0x21,
	0x2C, 0x03, 0x53, 0x06, 0x59, 0x28, 0x20, 0x3B, 0x7B, 0x36, 0x29, 0x0C,
	0x38, 0x05, 0x0E, 0x58, 0x2B, 0x1C, 0x37, 0x23, 0x0B, 0x18, 0x04, 0x11,
	0x18, 0x31, 0x01, 0x5D, 0x0B, 0x22, 0x59, 0x29, 0x5E, 0x06, 0x54, 0x23,
	0x0B, 0x39, 0x2B, 0x3D, 0x19, 0x5F, 0x5E, 0x01, 0x2A, 0x13, 0x39, 0x32,
	0x18, 0x36, 0x54, 0x5C, 0x02, 0x11, 0x43, 0x1B, 0x3B, 0x04, 0x0A, 0x39,
	0x16, 0x02, 0x1A, 0x36, 0x21, 0x33, 0x07, 0x0A, 0x71, 0x0D, 0x4E, 0x39,
	0x1E, 0x32, 0x0B, 0x25, 0x1C, 0x3D, 0x1B, 0x3F, 0x2C, 0x05, 0x0A, 0x7A,
	0x5D, 0x33, 0x22, 0x22, 0x3A, 0x2D, 0x3B, 0x5B, 0x32, 0x2B, 0x26, 0x1B,
	0x2F, 0x53, 0x28, 0x0F, 0x20, 0x1D, 0x02, 0x2C, 0x2D, 0x35, 0x05, 0x2E,
	0x3B, 0x25, 0x59, 0x2F, 0x40, 0x11, 0x39, 0x06, 0x04, 0x13, 0x03, 0x15,
	0x36, 0x38, 0x03, 0x07, 0x0A, 0x1B, 0x36, 0x23, 0x2E, 0x59, 0x0A, 0x5F,
	0x13, 0x7B, 0x35, 0x0D, 0x1A, 0x00, 0x6D, 0x5A, 0x04, 0x1E, 0x28, 0x32,
	0x2D, 0x17, 0x27, 0x40, 0x13, 0x2B, 0x55, 0x2A, 0x5E, 0x0E, 0x23, 0x20,
	0x26, 0x28, 0x0A, 0x07, 0x11, 0x3E, 0x0C, 0x15, 0x14, 0x55, 0x3B, 0x26,
	0x69, 0x38, 0x17, 0x38, 0x04, 0x09, 0x04, 0x31, 0x5F, 0x2E, 0x71, 0x55,
	0x0F, 0x34, 0x44, 0x12, 0x3F, 0x32, 0x23, 0x05, 0x05, 0x1A, 0x0A, 0x20,
	0x33, 0x70, 0x09, 0x2F, 0x45, 0x5A, 0x35, 0x34, 0x39, 0x0B, 0x1B, 0x38,
	0x1A, 0x33, 0x3D, 0x3A, 0x73, 0x1B, 0x2B, 0x3D, 0x22, 0x2F, 0x3F, 0x14,
	0x5E, 0x27, 0x11, 0x0E, 0x30, 0x21, 0x0A, 0x36, 0x00, 0x57, 0x34, 0x31,
	0x71, 0x2E, 0x13, 0x34, 0x28, 0x16, 0x27, 0x07, 0x1B, 0x01, 0x11, 0x18,
	0x2A, 0x25, 0x5D, 0x10, 0x19, 0x51, 0x26, 0x06, 0x0D, 0x58, 0x25, 0x56,
	0x2A, 0x32, 0x28, 0x29, 0x0A, 0x25, 0x12, 0x55, 0x08, 0x2C, 0x5C, 0x73,
	0x02, 0x26, 0x5B, 0x0D, 0x77, 0x01, 0x2B, 0x2F, 0x07, 0x25, 0x2E, 0x18,
	0x20, 0x38, 0x00, 0x22, 0x30, 0x29, 0x5E, 0x2B, 0x3E, 0x2C, 0x16, 0x5D,
	0x0A, 0x1B, 0x04, 0x34, 0x27, 0x3A, 0x25, 0x18, 0x27, 0x26, 0x20, 0x1C,
	0x15, 0x59, 0x1D, 0x16, 0x0A, 0x25, 0x57, 0x1F, 0x11, 0x43, 0x33, 0x36,
	0x2C, 0x75, 0x5E, 0x18, 0x5F, 0x32, 0x12, 0x08, 0x00, 0x0A, 0x39, 0x0B,
	0x25, 0x16, 0x45, 0x21, 0x09, 0x14, 0x07, 0x04, 0x03, 0x28, 0x1E, 0x34,
	0x5C, 0x52, 0x18, 0x1F, 0x50, 0x2A, 0x22, 0x1A, 0x34, 0x10, 0x0C, 0x52,
	0x75, 0x1E, 0x35, 0x38, 0x02, 0x35, 0x0B, 0x3B, 0x25, 0x40, 0x75, 0x1B,
	0x50, 0x34, 0x0D, 0x77, 0x08, 0x56, 0x04, 0x06, 0x31, 0x06, 0x33, 0x2A,
	0x1C, 0x0D, 0x04, 0x0F, 0x05, 0x25, 0x2E, 0x2B, 0x18, 0x2B, 0x2D, 0x3A,
	0x59, 0x07, 0x0B, 0x28, 0x38, 0x2E, 0x54, 0x2F, 0x5C, 0x30, 0x1E, 0x2C,
	0x57, 0x52, 0x0A, 0x19, 0x27, 0x14, 0x20, 0x29, 0x1F, 0x02, 0x5F, 0x5F,
	0x07, 0x5F, 0x38, 0x3B, 0x33, 0x0D, 0x0F, 0x0F, 0x06, 0x2F, 0x11, 0x38,
	0x14, 0x34, 0x27, 0x24, 0x3B, 0x2A, 0x18, 0x06, 0x3B, 0x43, 0x16, 0x28,
	0x3C, 0x28, 0x5F, 0x0B, 0x02, 0x38, 0x75, 0x3F, 0x0B, 0x28, 0x1F, 0x31,
	0x0D, 0x52, 0x05, 0x12, 0x0E, 0x5F, 0x4A, 0x02, 0x58, 0x69, 0x03, 0x2A,
	0x3F, 0x2D, 0x1B, 0x28, 0x34, 0x09, 0x23, 0x29, 0x16, 0x38, 0x2C, 0x08,
	0x6D, 0x04, 0x16, 0x08, 0x40, 0x27, 0x0B, 0x13, 0x5E, 0x5C, 0x70, 0x27,
	0x26, 0x1C, 0x00, 0x16, 0x3B, 0x17, 0x5E, 0x52, 0x0B, 0x08, 0x14, 0x3A,
	0x52, 0x3A, 0x15, 0x34, 0x5F, 0x20, 0x05, 0x1C, 0x54, 0x18, 0x3A, 0x2D,
	0x1D, 0x50, 0x1D, 0x24, 0x29, 0x5C, 0x19, 0x38, 0x01, 0x0E, 0x04, 0x4E,
	0x27, 0x59, 0x11, 0x3C, 0x51, 0x28, 0x2C, 0x2C, 0x14, 0x3B, 0x36, 0x21,
	0x07, 0x3D, 0x4E, 0x1C, 0x0C, 0x76, 0x3B, 0x0A, 0x41, 0x1B, 0x2B, 0x3B,
	0x2A, 0x0C, 0x11, 0x09, 0x00, 0x33, 0x05, 0x1A, 0x10, 0x08, 0x36, 0x19,
	0x05, 0x2E, 0x36, 0x30, 0x23, 0x3F, 0x1B, 0x2D, 0x18, 0x3A, 0x38, 0x34,
	0x0F, 0x00, 0x41, 0x53, 0x17, 0x07, 0x2D, 0x1B, 0x0D, 0x20, 0x20, 0x03,
	0x00, 0x13, 0x21, 0x38, 0x12, 0x18, 0x5F, 0x01, 0x55, 0x18, 0x00, 0x0E,
	0x09, 0x27, 0x56, 0x23, 0x44, 0x7B, 0x58, 0x2A, 0x17, 0x27, 0x31, 0x2D,
	0x14, 0x37, 0x3C, 0x10, 0x54, 0x32, 0x59, 0x12, 0x27, 0x36, 0x25, 0x5B,
	0x2C, 0x2B, 0x2D, 0x4E, 0x2C, 0x40, 0x10, 0x5F, 0x06, 0x2B, 0x12, 0x21,
	0x5A, 0x18, 0x3E, 0x0F, 0x25, 0x20, 0x16, 0x39, 0x00, 0x04, 0x59, 0x20,
	0x37, 0x00, 0x09, 0x23, 0x22, 0x0B, 0x44, 0x2F, 0x1A, 0x32, 0x2A, 0x11,
	0x09, 0x39, 0x25, 0x1B, 0x25, 0x17, 0x06, 0x57, 0x16, 0x19, 0x77, 0x2A,
	0x18, 0x24, 0x5E, 0x2C, 0x19, 0x2E, 0x41, 0x5E, 0x2A, 0x5F, 0x31, 0x3A,
	0x3B, 0x1A, 0x5C, 0x00, 0x21, 0x0A, 0x0C, 0x0E, 0x39, 0x34, 0x29, 0x27,
	0x59, 0x52, 0x29, 0x1D, 0x26, 0x1D, 0x4E, 0x0D, 0x0A, 0x36, 0x08, 0x25,
	0x5C, 0x5D, 0x04, 0x38, 0x0C, 0x3B, 0x06, 0x34, 0x5D, 0x0D, 0x2B, 0x58,
	0x77, 0x5C, 0x0D, 0x28, 0x20, 0x6D, 0x5A, 0x52, 0x2D, 0x1B, 0x06, 0x1B,
	0x50, 0x08, 0x5E, 0x7A, 0x21, 0x34, 0x3A, 0x22, 0x12, 0x1A, 0x26, 0x05,
	0x23, 0x3B, 0x2F, 0x0A, 0x00, 0x2D, 0x2A, 0x5A, 0x00, 0x1E, 0x32, 0x32,
	0x2A, 0x16, 0x1C, 0x11, 0x10, 0x27, 0x15, 0x57, 0x21, 0x0A, 0x22, 0x28,
	0x57, 0x22, 0x73, 0x5B, 0x06, 0x21, 0x1D, 0x13, 0x1D, 0x58, 0x3E, 0x3D,
	0x17, 0x03, 0x51, 0x0D, 0x21, 0x23, 0x3D, 0x0F, 0x59, 0x0D, 0x0C, 0x14,
	0x2F, 0x3F, 0x19, 0x01, 0x23, 0x11, 0x1A, 0x0A, 0x38, 0x03, 0x1B, 0x41,
	0x3C, 0x75, 0x5B, 0x25, 0x3C, 0x2A, 0x0F, 0x29, 0x30, 0x0C, 0x12, 0x04,
	0x0B, 0x4A, 0x5D, 0x01, 0x3A, 0x0E, 0x09, 0x5A, 0x5B, 0x37, 0x39, 0x4A,
	0x5F, 0x58, 0x0F, 0x2E, 0x14, 0x3C, 0x02, 0x13, 0x2E, 0x38, 0x3A, 0x18,
	0x07, 0x07, 0x4A, 0x58, 0x01, 0x32, 0x2F, 0x19, 0x5A, 0x07, 0x36, 0x39,
	0x22, 0x2C, 0x00, 0x2C, 0x0E, 0x2D, 0x37, 0x1F, 0x21, 0x26, 0x50, 0x5D,
	0x28, 0x3B, 0x3D, 0x38, 0x07, 0x1E, 0x08, 0x05, 0x31, 0x25, 0x0F, 0x30,
	0x3D, 0x2E, 0x04, 0x05, 0x70, 0x5A, 0x25, 0x38, 0x58, 0x1B, 0x2D, 0x02,
	0x2C, 0x0E, 0x16, 0x2E, 0x18, 0x19, 0x1D, 0x2F, 0x1A, 0x24, 0x04, 0x5C,
	0x32, 0x20, 0x59, 0x09, 0x31, 0x09, 0x26, 0x55, 0x56, 0x5F, 0x7B, 0x2D,
	0x10, 0x5C, 0x0E, 0x69, 0x14, 0x0A, 0x0D, 0x1E, 0x00, 0x5E, 0x32, 0x5B,
	0x3A, 0x06, 0x36, 0x27, 0x04, 0x31, 0x18, 0x0D, 0x19, 0x5B, 0x0E, 0x70,
	0x19, 0x11, 0x2A, 0x1B, 0x20, 0x38, 0x32, 0x1F, 0x59, 0x0D, 0x1F, 0x08,
	0x1B, 0x3B, 0x09, 0x5B, 0x22, 0x3A, 0x00, 0x33, 0x1E, 0x2B, 0x3A, 0x0F,
	0x30, 0x43, 0x29, 0x59, 0x59, 0x06, 0x59, 0x22, 0x57, 0x04, 0x2D, 0x59,
	0x54, 0x0D, 0x1F, 0x35, 0x02, 0x36, 0x21, 0x2A, 0x6D, 0x3C, 0x06, 0x5F,
	0x5D, 0x13, 0x02, 0x33, 0x29, 0x1D, 0x29, 0x38, 0x18, 0x2A, 0x13, 0x3A,
	0x02, 0x0E, 0x41, 0x53, 0x0C, 0x3F, 0x26, 0x26, 0x27, 0x2C, 0x2E, 0x56,
	0x5B, 0x02, 0x17, 0x0B, 0x59, 0x14, 0x1B, 0x01, 0x18, 0x0E, 0x1C, 0x5C,
	0x37, 0x3D, 0x54, 0x05, 0x3A, 0x29, 0x28, 0x00, 0x09, 0x2C, 0x35, 0x02,
	0x3B, 0x27, 0x40, 0x35, 0x1E, 0x26, 0x5A, 0x07, 0x77, 0x20, 0x25, 0x01,
	0x3B, 0x71, 0x08, 0x20, 0x1F, 0x44, 0x36, 0x35, 0x33, 0x18, 0x3F, 0x06,
	0x0A, 0x16, 0x39, 0x31, 0x17, 0x58, 0x23, 0x0D, 0x24, 0x08, 0x47, 0x4A,
	0x01, 0x1B, 0x25, 0x20, 0x0F, 0x04, 0x11, 0x24, 0x00, 0x52, 0x05, 0x1B,
	0x0B, 0x26, 0x02, 0x2C, 0x18, 0x2F, 0x26, 0x4A, 0x03, 0x03, 0x04, 0x18,
	0x0F, 0x06, 0x39, 0x29, 0x5F, 0x0A, 0x00, 0x22, 0x06, 0x01, 0x27, 0x34,
	0x0D, 0x21, 0x5B, 0x28, 0x1E, 0x24, 0x12, 0x5C, 0x32, 0x58, 0x22, 0x14,
	0x16, 0x35, 0x18, 0x1A, 0x0D, 0x3C, 0x33, 0x14, 0x12, 0x11, 0x0B, 0x28,
	0x06, 0x07, 0x2D, 0x04, 0x2E, 0x19, 0x32, 0x30, 0x29, 0x57, 0x3A, 0x38,
	0x2C, 0x39, 0x1B, 0x22, 0x2F, 0x36, 0x0A, 0x4E, 0x2F, 0x1D, 0x23, 0x0A,
	0x20, 0x3E, 0x22, 0x20, 0x3D, 0x22, 0x5B, 0x08, 0x13, 0x2B, 0x4A, 0x45,
	0x5F, 0x0A, 0x5B, 0x0D, 0x5B, 0x12, 0x71, 0x1B, 0x3B, 0x38, 0x5F, 0x36,
	0x29, 0x31, 0x24, 0x3F, 0x11, 0x1F, 0x50, 0x06, 0x3C, 0x3B, 0x3C, 0x33,
	0x04, 0x1A, 0x7B, 0x1E, 0x0E, 0x20, 0x3E, 0x12, 0x25, 0x2F, 0x0F, 0x5B,
	0x03, 0x3B, 0x35, 0x0B, 0x2F, 0x0F, 0x0B, 0x29, 0x2F, 0x27, 0x29, 0x08,
	0x0A, 0x23, 0x53, 0x01, 0x54, 0x0E, 0x45, 0x2A, 0x24, 0x26, 0x4A, 0x3F,
	0x23, 0x23, 0x26, 0x17, 0x41, 0x29, 0x08, 0x07, 0x29, 0x1C, 0x1D, 0x13,
	0x3E, 0x54, 0x5A, 0x28, 0x3B, 0x24, 0x2C, 0x2C, 0x06, 0x20, 0x5C, 0x16,
	0x5D, 0x3E, 0x69, 0x18, 0x0A, 0x36, 0x00, 0x25, 0x0F, 0x18, 0x5E, 0x03,
	0x08, 0x1B, 0x33, 0x59, 0x29, 0x15, 0x3D, 0x08, 0x3F, 0x20, 0x76, 0x24,
	0x09, 0x23, 0x44, 0x35, 0x07, 0x02, 0x04, 0x25, 0x0B, 0x3C, 0x2F, 0x34,
	0x3A, 0x30, 0x35, 0x4A, 0x17, 0x40, 0x1A, 0x5A, 0x2B, 0x1D, 0x03, 0x7A,
	0x08, 0x53, 0x29, 0x5D, 0x14, 0x54, 0x09, 0x37, 0x24, 0x76, 0x3F, 0x34,
	0x16, 0x38, 0x28, 0x58, 0x2D, 0x0C, 0x3A, 0x23, 0x1A, 0x59, 0x06, 0x23,
	0x1A, 0x0B, 0x09, 0x27, 0x2D, 0x3B, 0x2E, 0x2D, 0x2F, 0x0A, 0x29, 0x2E,
	0x12, 0x03, 0x5A, 0x10, 0x19, 0x17, 0x1F, 0x06, 0x29, 0x35, 0x4A, 0x2F,
	0x11, 0x04, 0x0F, 0x20, 0x45, 0x3A, 0x1B, 0x04, 0x59, 0x17, 0x5E, 0x72,
	0x22, 0x04, 0x3C, 0x3B, 0x13, 0x09, 0x00, 0x5D, 0x0C, 0x04, 0x15, 0x16,
	0x03, 0x24, 0x35, 0x14, 0x24, 0x38, 0x07, 0x74, 0x5E, 0x0C, 0x24, 0x0D,
	0x77, 0x1A, 0x0C, 0x2F, 0x33, 0x01, 0x0D, 0x30, 0x3B, 0x04, 0x0C, 0x5B,
	0x17, 0x2D, 0x40, 0x38, 0x29, 0x0D, 0x1C, 0x5A, 0x03, 0x5B, 0x28, 0x3A,
	0x00, 0x04, 0x1F, 0x23, 0x45, 0x38, 0x35, 0x0B, 0x39, 0x19, 0x23, 0x29,
	0x09, 0x16, 0x25, 0x1B, 0x10, 0x22, 0x39, 0x29, 0x3E, 0x0C, 0x0B, 0x18,
	0x57, 0x3C, 0x2C, 0x18, 0x26, 0x3E, 0x1C, 0x36, 0x18, 0x31, 0x01, 0x27,
	0x0B, 0x23, 0x2E, 0x18, 0x0C, 0x05, 0x0F, 0x0F, 0x34, 0x20, 0x15, 0x35,
	0x29, 0x34, 0x32, 0x13, 0x21, 0x0D, 0x02, 0x53, 0x2C, 0x0A, 0x36, 0x2B,
	0x08, 0x0D, 0x5E, 0x00, 0x38, 0x2C, 0x20, 0x1E, 0x27, 0x0B, 0x07, 0x27,
	0x3A, 0x55, 0x5D, 0x08, 0x01, 0x2A, 0x04, 0x45, 0x2D, 0x18, 0x2D, 0x17,
	0x2F, 0x23, 0x0B, 0x35, 0x0A, 0x2C, 0x53, 0x01, 0x0F, 0x0E, 0x0F, 0x3A,
	0x37, 0x3F, 0x2B, 0x07, 0x52, 0x36, 0x0B, 0x0D, 0x18, 0x18, 0x3B, 0x16,
	0x20, 0x26, 0x00, 0x2A, 0x25, 0x04, 0x1B, 0x38, 0x14, 0x02, 0x50, 0x06,
	0x04, 0x76, 0x43, 0x33, 0x21, 0x5F, 0x10, 0x5D, 0x59, 0x3D, 0x1B, 0x2D,
	0x18, 0x30, 0x25, 0x3A, 0x12, 0x07, 0x22, 0x29, 0x2A, 0x26, 0x07, 0x23,
	0x17, 0x2D, 0x74, 0x2E, 0x50, 0x27, 0x19, 0x14, 0x0D, 0x0E, 0x3E, 0x5B,
	0x69, 0x19, 0x35, 0x05, 0x0E, 0x70, 0x01, 0x05, 0x36, 0x00, 0x28, 0x1D,
	0x0F, 0x0B, 0x1B, 0x15, 0x2E, 0x51, 0x3D, 0x19, 0x2D, 0x22, 0x0D, 0x39,
	0x3F, 0x31, 0x04, 0x2B, 0x5A, 0x0E, 0x0C, 0x43, 0x26, 0x59, 0x03, 0x0D,
	0x2D, 0x0F, 0x24, 0x24, 0x1A, 0x01, 0x07, 0x06, 0x1A, 0x32, 0x5B, 0x06,
	0x17, 0x1B, 0x75, 0x2F, 0x54, 0x23, 0x38, 0x74, 0x3B, 0x2D, 0x27, 0x1C,
	0x74, 0x2F, 0x59, 0x28, 0x52, 0x21, 0x0D, 0x2F, 0x19, 0x18, 0x36, 0x47,
	0x59, 0x02, 0x27, 0x6D, 0x23, 0x11, 0x23, 0x29, 0x2F, 0x39, 0x03, 0x27,
	0x31, 0x05, 0x29, 0x37, 0x1C, 0x2A, 0x01, 0x36, 0x20, 0x3B, 0x2A, 0x70,
	0x2D, 0x52, 0x27, 0x52, 0x0B, 0x2E, 0x59, 0x29, 0x5E, 0x0F, 0x18, 0x2D,
	0x5E, 0x40, 0x32, 0x21, 0x50, 0x21, 0x0D, 0x30, 0x0F, 0x03, 0x24, 0x5B,
	0x77, 0x23, 0x06, 0x2B, 0x0A, 0x12, 0x3A, 0x0B, 0x3F, 0x29, 0x77, 0x09,
	0x0C, 0x1A, 0x31, 0x18, 0x5C, 0x12, 0x06, 0x01, 0x2E, 0x1A, 0x0A, 0x17,
	0x11, 0x35, 0x24, 0x0A, 0x16, 0x32, 0x00, 0x0F, 0x28, 0x1E, 0x2A, 0x25,
	0x5F, 0x23, 0x17, 0x3C, 0x00, 0x1C, 0x17, 0x24, 0x5D, 0x18, 0x00, 0x00,
	0x34, 0x0C, 0x05, 0x5C, 0x36, 0x09, 0x33, 0x0B, 0x09, 0x0A, 0x2F, 0x59,
	0x07, 0x02, 0x2A, 0x04, 0x53, 0x03, 0x20, 0x04, 0x3D, 0x08, 0x25, 0x23,
	0x38, 0x08, 0x44, 0x21, 0x2D, 0x10, 0x5C, 0x40, 0x03, 0x21, 0x0B, 0x36,
	0x2A, 0x24, 0x07, 0x2E, 0x27, 0x27, 0x7A, 0x01, 0x3B, 0x21, 0x06, 0x04,
	0x20, 0x15, 0x0A, 0x2D, 0x30, 0x15, 0x51, 0x3B, 0x11, 0x25, 0x1D, 0x14,
	0x28, 0x5C, 0x38, 0x3B, 0x29, 0x45, 0x40, 0x1A, 0x1A, 0x2F, 0x0F, 0x44,
	0x38, 0x0B, 0x11, 0x2F, 0x19, 0x25, 0x23, 0x0A, 0x2D, 0x18, 0x25, 0x5B,
	0x22, 0x28, 0x00, 0x29, 0x20, 0x2C, 0x0C, 0x58, 0x25, 0x54, 0x16, 0x41,
	0x2C, 0x01, 0x3F, 0x58, 0x19, 0x59, 0x7A, 0x3D, 0x2C, 0x05, 0x5C, 0x1B,
	0x39, 0x07, 0x56, 0x29, 0x30, 0x0A, 0x55, 0x2B, 0x12, 0x0E, 0x06, 0x39,
	0x45, 0x08, 0x2A, 0x16, 0x20, 0x36, 0x05, 0x18, 0x5A, 0x58, 0x24, 0x1A,
	0x2D, 0x04, 0x11, 0x34, 0x2F, 0x06, 0x26, 0x58, 0x09, 0x27, 0x35, 0x2A,
	0x0A, 0x3E, 0x08, 0x00, 0x0F, 0x15, 0x08, 0x19, 0x6D, 0x29, 0x0B, 0x21,
	0x1F, 0x72, 0x28, 0x0C, 0x3F, 0x3E, 0x00, 0x23, 0x20, 0x41, 0x20, 0x07,
	0x59, 0x35, 0x59, 0x12, 0x03, 0x07, 0x23, 0x03, 0x2A, 0x16, 0x27, 0x07,
	0x05, 0x23, 0x2C, 0x2F, 0x3B, 0x5F, 0x13, 0x0D, 0x3F, 0x27, 0x38, 0x53,
	0x77, 0x38, 0x05, 0x19, 0x20, 0x3A, 0x29, 0x58, 0x07, 0x24, 0x03, 0x5A,
	0x2F, 0x16, 0x28, 0x3B, 0x34, 0x2D, 0x3D, 0x5D, 0x06, 0x3B, 0x32, 0x45,
	0x39, 0x0F, 0x04, 0x36, 0x01, 0x31, 0x6D, 0x43, 0x23, 0x39, 0x3F, 0x0D,
	0x2D, 0x07, 0x25, 0x2E, 0x09, 0x47, 0x0A, 0x21, 0x13, 0x20, 0x16, 0x59,
	0x36, 0x2E, 0x0E, 0x2B, 0x08, 0x0C, 0x5D, 0x3A, 0x0B, 0x2B, 0x2A, 0x2F,
	0x77, 0x55, 0x18, 0x34, 0x0A, 0x0C, 0x5E, 0x37, 0x41, 0x05, 0x17, 0x2B,
	0x20, 0x0A, 0x00, 0x0D, 0x15, 0x2A, 0x0D, 0x29, 0x69, 0x3F, 0x0E, 0x06,
	0x39, 0x7A, 0x3E, 0x1B, 0x41, 0x38, 0x34, 0x25, 0x4E, 0x24, 0x12, 0x13,
	0x20, 0x0C, 0x2B, 0x01, 0x12, 0x39, 0x1B, 0x27, 0x28, 0x26, 0x24, 0x10,
	0x22, 0x52, 0x06, 0x1D, 0x0C, 0x3D, 0x1F, 0x7A, 0x59, 0x26, 0x24, 0x2A,
	0x14, 0x04, 0x2C, 0x17, 0x33, 0x34, 0x04, 0x57, 0x2F, 0x12, 0x06, 0x16,
	0x39, 0x05, 0x29, 0x37, 0x26, 0x00, 0x3F, 0x18, 0x75, 0x26, 0x59, 0x18,
	0x0C, 0x21, 0x15, 0x4E, 0x1C, 0x5B, 0x25, 0x1E, 0x0F, 0x5C, 0x01, 0x29,
	0x2A, 0x22, 0x28, 0x5C, 0x77, 0x38, 0x51, 0x3A, 0x18, 0x2E, 0x01, 0x16,
	0x3E, 0x44, 0x72, 0x1D, 0x4E, 0x14, 0x04, 0x34, 0x2D, 0x4A, 0x3F, 0x12,
	0x13, 0x26, 0x38, 0x3F, 0x08, 0x2E, 0x3E, 0x55, 0x5C, 0x3F, 0x72, 0x0B,
	0x34, 0x19, 0x20, 0x29, 0x2E, 0x02, 0x06, 0x24, 0x13, 0x2B, 0x55, 0x28,
	0x5E, 0x03, 0x59, 0x22, 0x57, 0x02, 0x26, 0x3B, 0x32, 0x00, 0x1D, 0x70,
	0x1E, 0x28, 0x14, 0x22, 0x77, 0x2A, 0x04, 0x06, 0x5A, 0x1A, 0x2A, 0x22,
	0x04, 0x04, 0x28, 0x47, 0x59, 0x5C, 0x1F, 0x01, 0x01, 0x0E, 0x03, 0x05,
	0x15, 0x35, 0x0C, 0x07, 0x31, 0x30, 0x29, 0x34, 0x03, 0x00, 0x30, 0x5B,
	0x58, 0x07, 0x06, 0x27, 0x1F, 0x05, 0x25, 0x52, 0x16, 0x04, 0x58, 0x16,
	0x5A, 0x11, 0x1C, 0x50, 0x26, 0x12, 0x2F, 0x5A, 0x2C, 0x5F, 0x2D, 0x36,
	0x3F, 0x58, 0x2A, 0x33, 0x01, 0x07, 0x2E, 0x3E, 0x0D, 0x21, 0x1C, 0x2A,
	0x41, 0x58, 0x76, 0x3B, 0x20, 0x18, 0x22, 0x05, 0x3D, 0x0D, 0x0F, 0x20,
	0x23, 0x2B, 0x24, 0x3A, 0x31, 0x0C, 0x58, 0x2B, 0x17, 0x22, 0x21, 0x2D,
	0x4A, 0x3A, 0x1F, 0x03, 0x1A, 0x06, 0x14, 0x22, 0x26, 0x47, 0x37, 0x14,
	0x52, 0x14, 0x34, 0x03, 0x5E, 0x3E, 0x00, 0x5A, 0x0F, 0x01, 0x1E, 0x15,
	0x47, 0x33, 0x00, 0x21, 0x7B, 0x2D, 0x09, 0x57, 0x40, 0x00, 0x09, 0x55,
	0x14, 0x07, 0x0C, 0x0A, 0x56, 0x17, 0x25, 0x16, 0x2D, 0x03, 0x05, 0x26,
	0x29, 0x27, 0x15, 0x0B, 0x05, 0x73, 0x0D, 0x54, 0x5F, 0x26, 0x2B, 0x0E,
	0x30, 0x25, 0x32, 0x0C, 0x15, 0x24, 0x5C, 0x2A, 0x24, 0x2E, 0x32, 0x3F,
	0x2A, 0x76, 0x28, 0x16, 0x3D, 0x33, 0x2D, 0x3F, 0x2E, 0x3F, 0x32, 0x3B,
	0x43, 0x16, 0x36, 0x22, 0x0D, 0x39, 0x22, 0x0B, 0x1D, 0x74, 0x1C, 0x30,
	0x07, 0x22, 0x14, 0x2B, 0x0C, 0x1C, 0x5C, 0x09, 0x00, 0x50, 0x02, 0x2A,
	0x01, 0x20, 0x4A, 0x07, 0x25, 0x07, 0x1E, 0x35, 0x2F, 0x11, 0x09, 0x55,
	0x06, 0x22, 0x3A, 0x03, 0x5E, 0x30, 0x00, 0x22, 0x20, 0x07, 0x20, 0x45,
	0x2F, 0x21, 0x04, 0x58, 0x06, 0x20, 0x3A, 0x3C, 0x4A, 0x00, 0x24, 0x7B,
	0x07, 0x33, 0x36, 0x03, 0x24, 0x2E, 0x23, 0x0F, 0x3B, 0x15, 0x0D, 0x50,
	0x04, 0x11, 0x35, 0x36, 0x0A, 0x21, 0x08, 0x16, 0x21, 0x10, 0x41, 0x0C,
	0x23, 0x03, 0x0F, 0x22, 0x28, 0x06, 0x07, 0x13, 0x57, 0x23, 0x35, 0x3C,
	0x15, 0x2F, 0x04, 0x08, 0x5A, 0x33, 0x22, 0x52, 0x08, 0x1B, 0x00, 0x34,
	0x2C, 0x35, 0x24, 0x54, 0x2B, 0x28, 0x00, 0x5F, 0x24, 0x1C, 0x21, 0x0B,
	0x0F, 0x29, 0x5C, 0x2F, 0x29, 0x24, 0x31, 0x2D, 0x53, 0x28, 0x15, 0x50,
	0x21, 0x01, 0x71, 0x3C, 0x50, 0x5A, 0x13, 0x37, 0x19, 0x2C, 0x5B, 0x01,
	0x27, 0x00, 0x19, 0x05, 0x3D, 0x14, 0x0B, 0x12, 0x36, 0x5A, 0x05, 0x1C,
	0x09, 0x04, 0x1F, 0x04, 0x3C, 0x52, 0x16, 0x20, 0x28, 0x55, 0x58, 0x1F,
	0x28, 0x2B, 0x2E, 0x0A, 0x3E, 0x03, 0x26, 0x5E, 0x1B, 0x1C, 0x38, 0x36,
	0x5E, 0x0F, 0x21, 0x5D, 0x0F, 0x01, 0x1B, 0x3C, 0x33, 0x2F, 0x0B, 0x50,
	0x3D, 0x26, 0x25, 0x19, 0x51, 0x36, 0x40, 0x37, 0x02, 0x14, 0x2A, 0x27,
	0x20, 0x25, 0x05, 0x39, 0x5C, 0x69, 0x55, 0x2B, 0x3A, 0x1C, 0x1B, 0x5F,
	0x31, 0x3B, 0x23, 0x0B, 0x2E, 0x28, 0x21, 0x3D, 0x27, 0x05, 0x37, 0x5C,
	0x00, 0x14, 0x2F, 0x0D, 0x3F, 0x5A, 0x1A, 0x1E, 0x59, 0x04, 0x1B, 0x71,
	0x39, 0x57, 0x1B, 0x5E, 0x25, 0x1A, 0x50, 0x45, 0x5F, 0x12, 0x03, 0x04,
	0x27, 0x28, 0x21, 0x2E, 0x04, 0x34, 0x02, 0x13, 0x25, 0x58, 0x22, 0x44,
	0x37, 0x18, 0x10, 0x36, 0x0E, 0x16, 0x58, 0x0B, 0x37, 0x01, 0x73, 0x00,
	0x20, 0x3D, 0x2D, 0x75, 0x07, 0x14, 0x57, 0x3D, 0x75, 0x22, 0x36, 0x3C,
	0x3E, 0x2C, 0x5D, 0x00, 0x00, 0x25, 0x15, 0x5C, 0x50, 0x56, 0x2D, 0x73,
	0x18, 0x06, 0x3E, 0x12, 0x12, 0x07, 0x2D, 0x03, 0x28, 0x24, 0x43, 0x51,
	0x17, 0x12, 0x06, 0x16, 0x2D, 0x5A, 0x29, 0x7A, 0x24, 0x54, 0x2C, 0x0D,
	0x03, 0x24, 0x2D, 0x2C, 0x25, 0x16, 0x5B, 0x18, 0x20, 0x2E, 0x06, 0x01,
	0x24, 0x04, 0x21, 0x06, 0x5A, 0x2E, 0x0B, 0x19, 0x2A, 0x29, 0x19, 0x0C,
	0x5E, 0x3B, 0x22, 0x54, 0x1C, 0x3E, 0x2D, 0x07, 0x02, 0x5F, 0x19, 0x0F,
	0x1F, 0x24, 0x20, 0x1C, 0x77, 0x34, 0x02, 0x0F, 0x21, 0x0A, 0x5E, 0x13,
	0x1A, 0x1C, 0x37, 0x36, 0x51, 0x05, 0x28, 0x36, 0x1B, 0x02, 0x00, 0x38,
	0x17, 0x5C, 0x37, 0x3E, 0x40, 0x03, 0x1C, 0x02, 0x5B, 0x5A, 0x37, 0x2D,
	0x4E, 0x2C, 0x28, 0x13, 0x1F, 0x55, 0x2D, 0x26, 0x1A, 0x09, 0x2F, 0x1C,
	0x19, 0x1B, 0x00, 0x13, 0x08, 0x21, 0x2F, 0x1C, 0x06, 0x22, 0x1C, 0x23,
	0x07, 0x26, 0x1D, 0x2A, 0x70, 0x3D, 0x35, 0x27, 0x3D, 0x2D, 0x29, 0x24,
	0x3F, 0x58, 0x70, 0x22, 0x3B, 0x02, 0x03, 0x12, 0x38, 0x08, 0x00, 0x3D,
	0x0F, 0x19, 0x4A, 0x2F, 0x3D, 0x2A, 0x54, 0x24, 0x5B, 0x2A, 0x37, 0x2D,
	0x07, 0x27, 0x24, 0x13, 0x24, 0x09, 0x28, 0x05, 0x69, 0x16, 0x56, 0x27,
	0x05, 0x03, 0x20, 0x0A, 0x04, 0x5F, 0x01, 0x21, 0x36, 0x17, 0x1D, 0x37,
	0x21, 0x22, 0x06, 0x33, 0x33, 0x5C, 0x29, 0x09, 0x12, 0x20, 0x14, 0x0E,
	0x1C, 0x0F, 0x6D, 0x1D, 0x27, 0x37, 0x29, 0x21, 0x28, 0x12, 0x07, 0x3D,
	0x25, 0x3C, 0x30, 0x2D, 0x3E, 0x2B, 0x3C, 0x0A, 0x36, 0x06, 0x04, 0x24,
	0x03, 0x3F, 0x0A, 0x18, 0x55, 0x16, 0x2C, 0x12, 0x00, 0x15, 0x23, 0x08,
	0x21, 0x2F, 0x3E, 0x59, 0x23, 0x03, 0x27, 0x5C, 0x3B, 0x56, 0x5C, 0x08,
	0x5A, 0x2B, 0x05, 0x05, 0x11, 0x09, 0x00, 0x09, 0x2C, 0x0F, 0x18, 0x4E,
	0x5B, 0x1E, 0x31, 0x25, 0x2E, 0x5D, 0x11, 0x09, 0x18, 0x07, 0x58, 0x3D,
	0x2E, 0x1B, 0x2E, 0x17, 0x29, 0x32, 0x2D, 0x23, 0x3F, 0x22, 0x1B, 0x25,
	0x26, 0x3D, 0x0D, 0x31, 0x59, 0x4A, 0x1D, 0x21, 0x0D, 0x3F, 0x35, 0x07,
	0x44, 0x0A, 0x19, 0x06, 0x5F, 0x0D, 0x7A, 0x2F, 0x54, 0x2B, 0x2D, 0x03,
	0x0A, 0x0A, 0x08, 0x22, 0x0A, 0x04, 0x26, 0x59, 0x0E, 0x0F, 0x1C, 0x50,
	0x18, 0x18, 0x35, 0x20, 0x22, 0x3C, 0x00, 0x30, 0x3C, 0x2A, 0x2C, 0x1E,
	0x13, 0x01, 0x00, 0x27, 0x3E, 0x1A, 0x07, 0x50, 0x1A, 0x24, 0x2D, 0x38,
	0x32, 0x20, 0x12, 0x0B, 0x38, 0x2B, 0x58, 0x3F, 0x09, 0x16, 0x2C, 0x1D,
	0x31, 0x03, 0x36, 0x13, 0x37, 0x38, 0x72, 0x27, 0x38, 0x5E, 0x44, 0x2F,
	0x2D, 0x52, 0x2A, 0x07, 0x34, 0x5E, 0x2F, 0x2B, 0x0A, 0x0E, 0x54, 0x17,
	0x2B, 0x27, 0x0E, 0x47, 0x30, 0x18, 0x08, 0x32, 0x43, 0x09, 0x02, 0x0A,
	0x0A, 0x3D, 0x31, 0x05, 0x5A, 0x2F, 0x0A, 0x54, 0x17, 0x26, 0x7B, 0x2D,
	0x54, 0x07, 0x1C, 0x25, 0x2A, 0x56, 0x58, 0x29, 0x3A, 0x1E, 0x17, 0x3F,
	0x11, 0x72, 0x55, 0x58, 0x09, 0x12, 0x6D, 0x16, 0x28, 0x05, 0x29, 0x27,
	0x3D, 0x02, 0x06, 0x5F, 0x2D, 0x34, 0x15, 0x08, 0x3A, 0x7A, 0x0B, 0x11,
	0x23, 0x0A, 0x27, 0x54, 0x27, 0x02, 0x19, 0x73, 0x29, 0x0F, 0x24, 0x32,
	0x3B, 0x22, 0x33, 0x2C, 0x31, 0x2A, 0x1F, 0x09, 0x0D, 0x40, 0x14, 0x1D,
	0x2A, 0x0D, 0x01, 0x21, 0x28, 0x12, 0x07, 0x52, 0x25, 0x24, 0x16, 0x0C,
	0x00, 0x12, 0x54, 0x20, 0x5B, 0x2A, 0x35, 0x0B, 0x54, 0x19, 0x29, 0x77,
	0x59, 0x13, 0x1F, 0x28, 0x77, 0x1B, 0x15, 0x3E, 0x22, 0x76, 0x38, 0x13,
	0x0B, 0x20, 0x11, 0x55, 0x3B, 0x0A, 0x2E, 0x74, 0x18, 0x19, 0x36, 0x05,
	0x14, 0x2A, 0x30, 0x0C, 0x44, 0x26, 0x59, 0x50, 0x38, 0x1A, 0x6D, 0x16,
	0x13, 0x57, 0x1C, 0x07, 0x59, 0x2C, 0x5C, 0x2A, 0x71, 0x29, 0x32, 0x27,
	0x58, 0x14, 0x22, 0x0B, 0x3C, 0x01, 0x24, 0x25, 0x29, 0x29, 0x3D, 0x07,
	0x55, 0x2E, 0x0D, 0x0D, 0x25, 0x1F, 0x19, 0x41, 0x2E, 0x75, 0x25, 0x4E,
	0x03, 0x0A, 0x73, 0x27, 0x2B, 0x1B, 0x1A, 0x76, 0x39, 0x4E, 0x3D, 0x5D,
	0x2B, 0x3B, 0x4E, 0x5E, 0x3C, 0x75, 0x5C, 0x22, 0x05, 0x28, 0x15, 0x2D,
	0x23, 0x27, 0x2A, 0x72, 0x2D, 0x39, 0x05, 0x3B, 0x0B, 0x26, 0x59, 0x2F,
	0x5E, 0x01, 0x2D, 0x09, 0x21, 0x53, 0x14, 0x54, 0x4A, 0x07, 0x2F, 0x0B,
	0x3C, 0x20, 0x16, 0x22, 0x76, 0x39, 0x51, 0x45, 0x53, 0x28, 0x3E, 0x20,
	0x36, 0x00, 0x28, 0x25, 0x07, 0x1F, 0x2D, 0x20, 0x2A, 0x0E, 0x22, 0x26,
	0x0C, 0x35, 0x30, 0x0D, 0x3C, 0x37, 0x34, 0x2A, 0x1C, 0x23, 0x7B, 0x38,
	0x14, 0x07, 0x25, 0x14, 0x25, 0x19, 0x1B, 0x0C, 0x73, 0x3A, 0x12, 0x27,
	0x06, 0x18, 0x14, 0x38, 0x04, 0x24, 0x33, 0x5B, 0x33, 0x59, 0x5C, 0x0F,
	0x19, 0x57, 0x2A, 0x3D, 0x2C, 0x35, 0x23, 0x56, 0x5F, 0x72, 0x5F, 0x53,
	0x36, 0x2A, 0x6D, 0x5B, 0x2D, 0x36, 0x5E, 0x0F, 0x15, 0x25, 0x3F, 0x13,
	0x17, 0x02, 0x56, 0x5F, 0x1B, 0x30, 0x38, 0x4A, 0x06, 0x1F, 0x0A, 0x3C,
	0x02, 0x24, 0x58, 0x3A, 0x0B, 0x38, 0x45, 0x53, 0x2A, 0x26, 0x22, 0x57,
	0x3A, 0x36, 0x22, 0x53, 0x09, 0x08, 0x3A, 0x15, 0x30, 0x20, 0x5F, 0x07,
	0x3F, 0x20, 0x14, 0x22, 0x70, 0x1B, 0x23, 0x5B, 0x23, 0x3B, 0x2F, 0x07,
	0x2F, 0x1E, 0x10, 0x47, 0x30, 0x05, 0x5D, 0x09, 0x1E, 0x4E, 0x16, 0x01,
	0x29, 0x3C, 0x0A, 0x02, 0x58, 0x71, 0x23, 0x00, 0x26, 0x3F, 0x0A, 0x39,
	0x22, 0x04, 0x00, 0x6D, 0x35, 0x00, 0x5C, 0x1C, 0x01, 0x1F, 0x00, 0x1D,
	0x0F, 0x73, 0x1F, 0x15, 0x39, 0x39, 0x2A, 0x1F, 0x00, 0x02, 0x0E, 0x72,
	0x1D, 0x0A, 0x5C, 0x1D, 0x0F, 0x59, 0x0D, 0x05, 0x21, 0x2D, 0x05, 0x59,
	0x1C, 0x59, 0x2F, 0x05, 0x50, 0x38, 0x28, 0x30, 0x29, 0x13, 0x20, 0x05,
	0x34, 0x00, 0x54, 0x0D, 0x1E, 0x17, 0x0A, 0x28, 0x56, 0x27, 0x69, 0x18,
	0x06, 0x22, 0x1C, 0x0A, 0x07, 0x2B, 0x1D, 0x21, 0x2F, 0x3F, 0x07, 0x58,
	0x59, 0x07, 0x2B, 0x30, 0x45, 0x38, 0x76, 0x0B, 0x11, 0x19, 0x2F, 0x77,
	0x21, 0x18, 0x28, 0x5C, 0x2A, 0x0A, 0x3B, 0x59, 0x38, 0x36, 0x2B, 0x39,
	0x03, 0x3D, 0x3A, 0x21, 0x57, 0x5D, 0x59, 0x18, 0x47, 0x30, 0x1A, 0x00,
	0x2E, 0x04, 0x2B, 0x17, 0x03, 0x75, 0x2D, 0x31, 0x38, 0x13, 0x05, 0x15,
	0x32, 0x41, 0x3A, 0x07, 0x16, 0x0C, 0x19, 0x53, 0x0B, 0x5B, 0x06, 0x07,
	0x3A, 0x2B, 0x0D, 0x2D, 0x1C, 0x44, 0x12, 0x2E, 0x0E, 0x06, 0x40, 0x30,
	0x43, 0x20, 0x24, 0x1C, 0x24, 0x3D, 0x2E, 0x3F, 0x5C, 0x35, 0x20, 0x18,
	0x5A, 0x59, 0x08, 0x0D, 0x56, 0x0A, 0x07, 0x21, 0x3B, 0x39, 0x04, 0x02,
	0x2E, 0x0D, 0x09, 0x0B, 0x1A, 0x10, 0x0E, 0x59, 0x38, 0x19, 0x69, 0x24,
	0x57, 0x5F, 0x11, 0x17, 0x5A, 0x18, 0x23, 0x1D, 0x0B, 0x23, 0x32, 0x3B,
	0x0E, 0x0B, 0x1C, 0x2D, 0x3F, 0x0A, 0x1B, 0x24, 0x0A, 0x3E, 0x3E, 0x01,
	0x58, 0x3B, 0x29, 0x19, 0x16, 0x29, 0x59, 0x06, 0x26, 0x35, 0x05, 0x15,
	0x0C, 0x06, 0x20, 0x07, 0x59, 0x3F, 0x33, 0x2C, 0x27, 0x30, 0x58, 0x29,
	0x38, 0x20, 0x59, 0x2D, 0x53, 0x2B, 0x2D, 0x09, 0x1B, 0x53, 0x15, 0x0E,
	0x31, 0x19, 0x26, 0x3B, 0x06, 0x16, 0x2A, 0x12, 0x75, 0x26, 0x2A, 0x3E,
	0x1D, 0x0B, 0x05, 0x30, 0x01, 0x5B, 0x29, 0x0A, 0x57, 0x56, 0x1E, 0x0F,
	0x08, 0x29, 0x28, 0x2D, 0x0C, 0x58, 0x0A, 0x1D, 0x03, 0x0D, 0x19, 0x16,
	0x5B, 0x02, 0x69, 0x25, 0x13, 0x41, 0x12, 0x71, 0x3D, 0x08, 0x0C, 0x0C,
	0x24, 0x36, 0x13, 0x5F, 0x39, 0x37, 0x2A, 0x26, 0x5E, 0x33, 0x7B, 0x5E,
	0x16, 0x36, 0x33, 0x70, 0x2D, 0x39, 0x27, 0x32, 0x29, 0x2E, 0x2E, 0x2F,
	0x44, 0x00, 0x0D, 0x30, 0x24, 0x5E, 0x14, 0x55, 0x54, 0x26, 0x06, 0x03,
	0x1A, 0x2A, 0x17, 0x08, 0x14, 0x1F, 0x16, 0x5C, 0x0D, 0x10, 0x59, 0x0A,
	0x1C, 0x02, 0x16, 0x07, 0x02, 0x3E, 0x20, 0x27, 0x09, 0x35, 0x45, 0x22,
	0x28, 0x21, 0x39, 0x16, 0x1D, 0x69, 0x18, 0x28, 0x1E, 0x1D, 0x36, 0x2F,
	0x50, 0x59, 0x27, 0x23, 0x2D, 0x15, 0x0B, 0x5E, 0x01, 0x36, 0x25, 0x0A,
	0x0C, 0x0C, 0x15, 0x07, 0x59, 0x2D, 0x1B, 0x00, 0x0B, 0x36, 0x5B, 0x00,
	0x1A, 0x52, 0x3A, 0x08, 0x21, 0x0A, 0x0F, 0x18, 0x5B, 0x0D, 0x03, 0x51,
	0x27, 0x23, 0x7A, 0x2E, 0x3B, 0x26, 0x27, 0x2D, 0x25, 0x1B, 0x23, 0x29,
	0x2F, 0x39, 0x17, 0x27, 0x02, 0x27, 0x3E, 0x2B, 0x38, 0x5A, 0x24, 0x28,
	0x12, 0x28, 0x07, 0x0B, 0x16, 0x57, 0x5D, 0x3A, 0x0F, 0x1D, 0x4A, 0x2A,
	0x3D, 0x2A, 0x15, 0x26, 0x5D, 0x28, 0x20, 0x1F, 0x4A, 0x3B, 0x2C, 0x13,
	0x5E, 0x32, 0x29, 0x3A, 0x2D, 0x22, 0x32, 0x01, 0x00, 0x23, 0x54, 0x3B,
	0x26, 0x03, 0x15, 0x3E, 0x51, 0x01, 0x52, 0x00, 0x1D, 0x59, 0x56, 0x2F,
	0x7A, 0x07, 0x50, 0x2F, 0x1D, 0x2B, 0x09, 0x30, 0x0D, 0x01, 0x14, 0x1E,
	0x19, 0x24, 0x5B, 0x2B, 0x01, 0x00, 0x5F, 0x02, 0x0E, 0x3C, 0x59, 0x2C,
	0x19, 0x28, 0x23, 0x14, 0x04, 0x11, 0x11, 0x07, 0x08, 0x2D, 0x3B, 0x26,
	0x28, 0x54, 0x29, 0x3F, 0x34, 0x47, 0x57, 0x2A, 0x0F, 0x7A, 0x05, 0x28,
	0x5C, 0x0D, 0x2E, 0x20, 0x1B, 0x57, 0x3C, 0x0D, 0x27, 0x56, 0x38, 0x1C,
	0x16, 0x18, 0x05, 0x2B, 0x04, 0x24, 0x07, 0x17, 0x28, 0x5D, 0x71, 0x5A,
	0x0E, 0x04, 0x2F, 0x29, 0x38, 0x34, 0x05, 0x05, 0x2A, 0x0F, 0x1B, 0x1C,
	0x38, 0x05, 0x36, 0x07, 0x19, 0x07, 0x75, 0x26, 0x58, 0x25, 0x3F, 0x27,
	0x3F, 0x25, 0x24, 0x23, 0x3A, 0x24, 0x0B, 0x08, 0x3A, 0x0F, 0x0B, 0x3B,
	0x5A, 0x3D, 0x36, 0x08, 0x25, 0x5D, 0x0E, 0x76, 0x2E, 0x54, 0x2A, 0x52,
	0x25, 0x2E, 0x16, 0x2D, 0x5E, 0x03, 0x0B, 0x09, 0x3E, 0x32, 0x0E, 0x1E,
	0x4A, 0x5A, 0x3A, 0x21, 0x29, 0x0F, 0x0C, 0x27, 0x38, 0x5A, 0x29, 0x38,
	0x1C, 0x76, 0x2D, 0x59, 0x1A, 0x1F, 0x7B, 0x24, 0x0F, 0x05, 0x58, 0x0B,
	0x38, 0x13, 0x26, 0x12, 0x69, 0x2B, 0x10, 0x3F, 0x1E, 0x10, 0x02, 0x04,
	0x08, 0x2A, 0x6D, 0x25, 0x50, 0x2F, 0x28, 0x77, 0x0B, 0x3B, 0x2C, 0x5A,
	0x35, 0x1E, 0x03, 0x5B, 0x26, 0x0F, 0x04, 0x59, 0x29, 0x1B, 0x03, 0x1A,
	0x20, 0x41, 0x22, 0x34, 0x0B, 0x29, 0x17, 0x44, 0x12, 0x5A, 0x51, 0x25,
	0x38, 0x04, 0x55, 0x3B, 0x1E, 0x1C, 0x72, 0x3B, 0x19, 0x01, 0x04, 0x34,
	0x09, 0x23, 0x1E, 0x0A, 0x6D, 0x36, 0x26, 0x3F, 0x3A, 0x76, 0x02, 0x52,
	0x16, 0x58, 0x33, 0x5D, 0x53, 0x2C, 0x1F, 0x77, 0x21, 0x0A, 0x56, 0x31,
	0x0B, 0x2E, 0x51, 0x1A, 0x0E, 0x37, 0x0E, 0x27, 0x06, 0x24, 0x35, 0x39,
	0x0E, 0x58, 0x00, 0x70, 0x07, 0x27, 0x37, 0x25, 0x0F, 0x02, 0x11, 0x5F,
	0x1C, 0x0D, 0x0A, 0x00, 0x16, 0x0A, 0x70, 0x29, 0x15, 0x5D, 0x3E, 0x24,
	0x25, 0x03, 0x0F, 0x3C, 0x2A, 0x39, 0x00, 0x21, 0x02, 0x73, 0x36, 0x0A,
	0x5C, 0x59, 0x11, 0x1F, 0x28, 0x3E, 0x1C, 0x09, 0x1E, 0x0F, 0x16, 0x03,
	0x3A, 0x39, 0x04, 0x0B, 0x33, 0x07, 0x01, 0x13, 0x2B, 0x21, 0x36, 0x14,
	0x20, 0x3A, 0x21, 0x38, 0x2D, 0x03, 0x05, 0x38, 0x29, 0x2D, 0x0E, 0x06,
	0x21, 0x77, 0x23, 0x12, 0x04, 0x12, 0x06, 0x35, 0x39, 0x21, 0x2E, 0x7B,
	0x58, 0x27, 0x23, 0x27, 0x20, 0x03, 0x18, 0x01, 0x2F, 0x23, 0x5D, 0x53,
	0x3E, 0x26, 0x2E, 0x24, 0x52, 0x09, 0x2E, 0x3B, 0x24, 0x18, 0x38, 0x00,
	0x2E, 0x47, 0x09, 0x04, 0x40, 0x35, 0x0B, 0x54, 0x38, 0x29, 0x06, 0x59,
	0x17, 0x0A, 0x2F, 0x33, 0x22, 0x22, 0x2C, 0x3B, 0x70, 0x07, 0x23, 0x0B,
	0x00, 0x34, 0x0B, 0x57, 0x05, 0x11, 0x20, 0x58, 0x2C, 0x02, 0x26, 0x00,
	0x19, 0x36, 0x3C, 0x2F, 0x15, 0x04, 0x05, 0x0A, 0x22, 0x35, 0x18, 0x20,
	0x34, 0x0C, 0x17, 0x0B, 0x20, 0x5A, 0x2F, 0x21, 0x3D, 0x2C, 0x06, 0x0E,
	0x07, 0x34, 0x4E, 0x45, 0x5F, 0x0B, 0x0D, 0x51, 0x3B, 0x1B, 0x7B, 0x2B,
	0x03, 0x01, 0x0F, 0x15, 0x55, 0x16, 0x2A, 0x12, 0x13, 0x5C, 0x2D, 0x21,
	0x28, 0x30, 0x43, 0x18, 0x20, 0x13, 0x34, 0x54, 0x52, 0x20, 0x3F, 0x0A,
	0x0E, 0x2F, 0x3D, 0x39, 0x05, 0x05, 0x02, 0x03, 0x18, 0x7B, 0x2B, 0x4E,
	0x14, 0x05, 0x3A, 0x2D, 0x50, 0x09, 0x27, 0x11, 0x2D, 0x26, 0x3F, 0x23,
	0x0B, 0x28, 0x02, 0x22, 0x03, 0x12, 0x3E, 0x02, 0x3B, 0x20, 0x2C, 0x24,
	0x35, 0x3D, 0x07, 0x38, 0x26, 0x56, 0x3A, 0x5D, 0x09, 0x05, 0x25, 0x41,
	0x2F, 0x31, 0x05, 0x17, 0x2F, 0x0D, 0x2C, 0x06, 0x33, 0x1A, 0x59, 0x28,
	0x5C, 0x08, 0x41, 0x5F, 0x75, 0x27, 0x0E, 0x1C, 0x1C, 0x3A, 0x36, 0x00,
	0x1B, 0x0E, 0x08, 0x1D, 0x53, 0x04, 0x5D, 0x73, 0x2A, 0x55, 0x58, 0x5B,
	0x32, 0x2E, 0x0B, 0x0A, 0x27, 0x74, 0x16, 0x57, 0x38, 0x5C, 0x76, 0x21,
	0x0A, 0x2D, 0x3C, 0x03, 0x1E, 0x20, 0x39, 0x1E, 0x2D, 0x3B, 0x2D, 0x28,
	0x53, 0x3B, 0x35, 0x53, 0x05, 0x00, 0x3B, 0x34, 0x50, 0x21, 0x2D, 0x35,
	0x02, 0x30, 0x56, 0x2A, 0x21, 0x1E, 0x15, 0x2F, 0x0E, 0x0C, 0x0D, 0x2D,
	0x06, 0x06, 0x37, 0x09, 0x1B, 0x24, 0x0F, 0x08, 0x59, 0x13, 0x07, 0x22,
	0x7A, 0x02, 0x51, 0x0A, 0x19, 0x2C, 0x23, 0x02, 0x05, 0x3B, 0x04, 0x2F,
	0x03, 0x41, 0x1C, 0x0D, 0x36, 0x20, 0x1F, 0x5A, 0x36, 0x2F, 0x2A, 0x1C,
	0x39, 0x32, 0x58, 0x2E, 0x21, 0x11, 0x36, 0x01, 0x20, 0x22, 0x20, 0x17,
	0x07, 0x2B, 0x5D, 0x28, 0x21, 0x5E, 0x0A, 0x3F, 0x08, 0x2E, 0x2F, 0x2C,
	0x1E, 0x05, 0x26, 0x2E, 0x10, 0x5F, 0x59, 0x03, 0x0A, 0x2B, 0x17, 0x3A,
	0x27, 0x3D, 0x37, 0x5D, 0x2D, 0x0C, 0x14, 0x27, 0x3D, 0x21, 0x24, 0x3D,
	0x59, 0x41, 0x0F, 0x03, 0x1D, 0x4A, 0x56, 0x28, 0x21, 0x04, 0x2A, 0x3F,
	0x58, 0x3A, 0x2E, 0x18, 0x25, 0x27, 0x04, 0x2D, 0x0E, 0x05, 0x1B, 0x6D,
	0x1A, 0x37, 0x06, 0x25, 0x16, 0x15, 0x39, 0x39, 0x26, 0x2C, 0x54, 0x36,
	0x1C, 0x3D, 0x32, 0x04, 0x34, 0x0A, 0x07, 0x14, 0x1C, 0x55, 0x3B, 0x2D,
	0x69, 0x5B, 0x32, 0x58, 0x0D, 0x69, 0x39, 0x39, 0x2B, 0x33, 0x0E, 0x16,
	0x35, 0x28, 0x0D, 0x2F, 0x07, 0x13, 0x1C, 0x1E, 0x2A, 0x47, 0x0A, 0x37,
	0x33, 0x07, 0x34, 0x28, 0x3B, 0x31, 0x0A, 0x16, 0x19, 0x05, 0x1E, 0x69,
	0x1C, 0x55, 0x36, 0x0E, 0x2B, 0x21, 0x53, 0x38, 0x5B, 0x71, 0x24, 0x57,
	0x0A, 0x00, 0x08, 0x01, 0x39, 0x21, 0x02, 0x69, 0x06, 0x30, 0x56, 0x3A,
	0x31, 0x00, 0x53, 0x1D, 0x1F, 0x2C, 0x47, 0x02, 0x05, 0x2C, 0x71, 0x2F,
	0x25, 0x18, 0x53, 0x05, 0x25, 0x38, 0x0A, 0x2D, 0x0A, 0x5F, 0x14, 0x19,
	0x05, 0x32, 0x59, 0x32, 0x0F, 0x01, 0x13, 0x07, 0x13, 0x29, 0x2F, 0x69,
	0x18, 0x52, 0x09, 0x1E, 0x2F, 0x05, 0x4A, 0x07, 0x12, 0x2A, 0x36, 0x4E,
	0x18, 0x05, 0x2A, 0x1F, 0x16, 0x5C, 0x52, 0x73, 0x2B, 0x32, 0x28, 0x23,
	0x00, 0x0A, 0x12, 0x0C, 0x3A, 0x09, 0x35, 0x2A, 0x17, 0x27, 0x00, 0x2D,
	0x2A, 0x02, 0x2C, 0x75, 0x5E, 0x30, 0x16, 0x09, 0x77, 0x07, 0x35, 0x5A,
	0x12, 0x15, 0x0E, 0x12, 0x57, 0x29, 0x23, 0x06, 0x2C, 0x24, 0x3E, 0x2A,
	0x1A, 0x37, 0x2B, 0x1D, 0x73, 0x36, 0x13, 0x03, 0x27, 0x05, 0x3C, 0x03,
	0x19, 0x52, 0x7A, 0x20, 0x37, 0x41, 0x5D, 0x1B, 0x3D, 0x28, 0x25, 0x03,
	0x72, 0x0B, 0x22, 0x3E, 0x52, 0x74, 0x00, 0x08, 0x0A, 0x3B, 0x7A, 0x55,
	0x15, 0x26, 0x04, 0x03, 0x07, 0x2E, 0x56, 0x2A, 0x21, 0x04, 0x10, 0x3F,
	0x44, 0x35, 0x3C, 0x28, 0x03, 0x20, 0x23, 0x3C, 0x31, 0x2C, 0x3C, 0x13,
	0x59, 0x19, 0x25, 0x12, 0x1A, 0x54, 0x1B, 0x5A, 0x08, 0x35, 0x00, 0x3B,
	0x22, 0x06, 0x38, 0x3E, 0x50, 0x16, 0x24, 0x3B, 0x3F, 0x18, 0x2F, 0x2F,
	0x38, 0x0E, 0x33, 0x0F, 0x19, 0x75, 0x29, 0x2A, 0x5A, 0x26, 0x2D, 0x0A,
	0x2B, 0x39, 0x38, 0x71, 0x47, 0x2E, 0x58, 0x0D, 0x00, 0x59, 0x0C, 0x2A,
	0x0C, 0x00, 0x1B, 0x27, 0x5B, 0x26, 0x05, 0x01, 0x03, 0x41, 0x1D, 0x7B,
	0x22, 0x18, 0x28, 0x05, 0x3A, 0x3A, 0x08, 0x45, 0x08, 0x00, 0x23, 0x2F,
	0x3D, 0x1F, 0x07, 0x3C, 0x2B, 0x5C, 0x13, 0x09, 0x0D, 0x57, 0x1A, 0x1A,
	0x77, 0x24, 0x0C, 0x2B, 0x19, 0x00, 0x09, 0x1B, 0x14, 0x24, 0x15, 0x0E,
	0x07, 0x25, 0x5E, 0x14, 0x0B, 0x2D, 0x3F, 0x59, 0x32, 0x0A, 0x39, 0x00,
	0x11, 0x18, 0x1B, 0x22, 0x23, 0x05, 0x21, 0x2E, 0x59, 0x06, 0x3D, 0x03,
	0x0A, 0x06, 0x14, 0x22, 0x0E, 0x1B, 0x25, 0x5B, 0x2A, 0x3B, 0x2E, 0x31,
	0x1E, 0x5C, 0x2C, 0x0B, 0x0C, 0x22, 0x28, 0x07, 0x26, 0x19, 0x20, 0x38,
	0x04, 0x08, 0x58, 0x07, 0x25, 0x37, 0x38, 0x26, 0x36, 0x1C, 0x77, 0x25,
	0x25, 0x17, 0x28, 0x20, 0x2D, 0x2F, 0x05, 0x2C, 0x3B, 0x20, 0x15, 0x5B,
	0x21, 0x2A, 0x20, 0x57, 0x45, 0x33, 0x0F, 0x0B, 0x59, 0x19, 0x5A, 0x03,
	0x0A, 0x06, 0x3A, 0x22, 0x05, 0x39, 0x20, 0x0B, 0x29, 0x3A, 0x24, 0x27,
	0x1E, 0x1C, 0x2F, 0x29, 0x05, 0x24, 0x5B, 0x09, 0x59, 0x11, 0x5A, 0x3C,
	0x76, 0x5E, 0x12, 0x58, 0x1F, 0x0A, 0x03, 0x50, 0x27, 0x2D, 0x26, 0x24,
	0x00, 0x0A, 0x3D, 0x74, 0x5C, 0x50, 0x0D, 0x21, 0x27, 0x09, 0x09, 0x1F,
	0x52, 0x3B, 0x02, 0x04, 0x2D, 0x0A, 0x71, 0x5E, 0x20, 0x22, 0x22, 0x12,
	0x07, 0x22, 0x56, 0x28, 0x7A, 0x05, 0x50, 0x2F, 0x0D, 0x25, 0x02, 0x28,
	0x23, 0x59, 0x0B, 0x0A, 0x0C, 0x3F, 0x09, 0x0B, 0x0D, 0x16, 0x2D, 0x5E,
	0x01, 0x1C, 0x20, 0x0B, 0x59, 0x01, 0x5D, 0x38, 0x27, 0x1B, 0x2F, 0x06,
	0x0E, 0x04, 0x52, 0x34, 0x26, 0x53, 0x3D, 0x33, 0x05, 0x24, 0x26, 0x5D,
	0x1C, 0x2C, 0x39, 0x4A, 0x2D, 0x53, 0x28, 0x34, 0x20, 0x08, 0x00, 0x12,
	0x3D, 0x29, 0x5A, 0x25, 0x3B, 0x26, 0x31, 0x0C, 0x31, 0x0B, 0x47, 0x2A,
	0x08, 0x01, 0x2B, 0x18, 0x56, 0x0D, 0x18, 0x31, 0x2E, 0x14, 0x3C, 0x0A,
	0x13, 0x26, 0x10, 0x2F, 0x44, 0x03, 0x5C, 0x06, 0x1B, 0x1C, 0x06, 0x59,
	0x2B, 0x2D, 0x23, 0x0C, 0x36, 0x20, 0x39, 0x29, 0x18, 0x03, 0x05, 0x17,
	0x1E, 0x7B, 0x0E, 0x51, 0x00, 0x1C, 0x36, 0x0D, 0x0F, 0x3F, 0x27, 0x29,
	0x5D, 0x55, 0x2A, 0x53, 0x2A, 0x36, 0x23, 0x1A, 0x1C, 0x37, 0x5A, 0x05,
	0x3E, 0x24, 0x28, 0x20, 0x17, 0x2C, 0x12, 0x13, 0x23, 0x38, 0x2D, 0x18,
	0x03, 0x23, 0x32, 0x20, 0x0C, 0x0F, 0x3F, 0x20, 0x18, 0x29, 0x27, 0x3D,
	0x0B, 0x19, 0x2D, 0x3B, 0x26, 0x18, 0x2C, 0x0D, 0x0B, 0x47, 0x32, 0x27,
	0x40, 0x00, 0x35, 0x4E, 0x2F, 0x1B, 0x29, 0x20, 0x09, 0x02, 0x12, 0x29,
	0x18, 0x08, 0x3B, 0x04, 0x36, 0x39, 0x10, 0x14, 0x31, 0x72, 0x01, 0x3B,
	0x07, 0x5D, 0x14, 0x21, 0x36, 0x21, 0x26, 0x32, 0x16, 0x11, 0x17, 0x24,
	0x20, 0x0F, 0x07, 0x09, 0x5F, 0x2B, 0x24, 0x4E, 0x17, 0x1A, 0x31, 0x2D,
	0x53, 0x3F, 0x01, 0x0B, 0x36, 0x0A, 0x2A, 0x0E, 0x03, 0x0F, 0x06, 0x0B,
	0x3A, 0x0D, 0x58, 0x25, 0x5B, 0x2D, 0x7A, 0x29, 0x51, 0x02, 0x0D, 0x15,
	0x5C, 0x3B, 0x34, 0x1F, 0x35, 0x05, 0x2D, 0x58, 0x2F, 0x3B, 0x24, 0x35,
	0x14, 0x1A, 0x38, 0x2D, 0x59, 0x5C, 0x0E, 0x76, 0x54, 0x09, 0x23, 0x58,
	0x74, 0x5D, 0x31, 0x0F, 0x52, 0x16, 0x1F, 0x2C, 0x00, 0x32, 0x0B, 0x5B,
	0x10, 0x0D, 0x1C, 0x29, 0x19, 0x2C, 0x5A, 0x18, 0x13, 0x23, 0x38, 0x2C,
	0x08, 0x37, 0x5D, 0x0C, 0x08, 0x31, 0x18, 0x5A, 0x4A, 0x00, 0x33, 0x74,
	0x2F, 0x2F, 0x05, 0x1A, 0x29, 0x2E, 0x09, 0x0F, 0x1D, 0x10, 0x19, 0x30,
	0x5C, 0x1C, 0x01, 0x59, 0x22, 0x5B, 0x29, 0x6D, 0x25, 0x14, 0x3D, 0x04,
	0x3B, 0x2B, 0x35, 0x45, 0x1F, 0x32, 0x2D, 0x3B, 0x1A, 0x29, 0x7B, 0x3A,
	0x15, 0x3E, 0x1B, 0x12, 0x19, 0x2C, 0x5B, 0x1D, 0x03, 0x24, 0x0F, 0x29,
	0x18, 0x0B, 0x55, 0x51, 0x2D, 0x38, 0x10, 0x19, 0x33, 0x25, 0x31, 0x2B,
	0x05, 0x22, 0x1B, 0x11, 0x07, 0x00, 0x0E, 0x5F, 0x28, 0x06, 0x07, 0x10,
	0x5B, 0x1B, 0x13, 0x3C, 0x06, 0x23, 0x13, 0x27, 0x3D, 0x25, 0x5B, 0x23,
	0x3B, 0x24, 0x03, 0x16, 0x13, 0x25, 0x58, 0x32, 0x23, 0x07, 0x2E, 0x35,
	0x23, 0x0A, 0x40, 0x03, 0x3A, 0x0B, 0x56, 0x28, 0x18, 0x2F, 0x31, 0x37,
	0x06, 0x24, 0x54, 0x27, 0x23, 0x06, 0x0D, 0x5E, 0x00, 0x21, 0x3F, 0x01,
	0x59, 0x2C, 0x1C, 0x3B, 0x71, 0x09, 0x2D, 0x22, 0x33, 0x07, 0x1E, 0x28,
	0x0B, 0x06, 0x07, 0x5D, 0x39, 0x3B, 0x3B, 0x0B, 0x2D, 0x59, 0x25, 0x06,
	0x71, 0x3D, 0x08, 0x1A, 0x09, 0x2B, 0x3E, 0x0A, 0x00, 0x25, 0x06, 0x3C,
	0x0F, 0x19, 0x20, 0x18, 0x1E, 0x16, 0x22, 0x12, 0x75, 0x58, 0x25, 0x56,
	0x23, 0x32, 0x2D, 0x0F, 0x18, 0x1F, 0x2E, 0x24, 0x39, 0x18, 0x19, 0x2F,
	0x55, 0x20, 0x3C, 0x38, 0x2D, 0x5A, 0x2C, 0x27, 0x3C, 0x11, 0x09, 0x12,
	0x1E, 0x02, 0x37, 0x0B, 0x50, 0x0C, 0x3C, 0x03, 0x0E, 0x20, 0x26, 0x00,
	0x20, 0x35, 0x32, 0x0D, 0x2D, 0x26, 0x1E, 0x0C, 0x3F, 0x5F, 0x16, 0x1F,
	0x26, 0x0B, 0x0D, 0x33, 0x16, 0x2D, 0x1D, 0x31, 0x11, 0x08, 0x54, 0x3E,
	0x05, 0x71, 0x2A, 0x05, 0x26, 0x03, 0x00, 0x5E, 0x56, 0x41, 0x0D, 0x25,
	0x15, 0x0B, 0x56, 0x2D, 0x77, 0x2F, 0x58, 0x18, 0x5A, 0x37, 0x27, 0x2E,
	0x00, 0x09, 0x06, 0x3A, 0x0D, 0x5D, 0x00, 0x77, 0x25, 0x29, 0x21, 0x58,
	0x32, 0x05, 0x07, 0x22, 0x06, 0x3B, 0x0F, 0x0D, 0x5B, 0x22, 0x04, 0x07,
	0x39, 0x3E, 0x39, 0x2E, 0x36, 0x0B, 0x2B, 0x3D, 0x76, 0x38, 0x11, 0x1A,
	0x3A, 0x31, 0x0D, 0x2D, 0x1C, 0x58, 0x35, 0x1E, 0x18, 0x26, 0x1C, 0x15,
	0x07, 0x2A, 0x56, 0x3F, 0x21, 0x07, 0x11, 0x56, 0x5E, 0x18, 0x47, 0x23,
	0x14, 0x2E, 0x14, 0x1A, 0x02, 0x3C, 0x2E, 0x23, 0x00, 0x2E, 0x3B, 0x59,
	0x15, 0x19, 0x3B, 0x18, 0x53, 0x18, 0x29, 0x3B, 0x06, 0x26, 0x35, 0x38,
	0x52, 0x1D, 0x58, 0x30, 0x3D, 0x04, 0x37, 0x38, 0x3B, 0x26, 0x05, 0x37,
	0x29, 0x38, 0x27, 0x50, 0x1A, 0x5D, 0x11, 0x3A, 0x06, 0x3A, 0x3E, 0x3B,
	0x43, 0x2B, 0x0C, 0x5B, 0x26, 0x2B, 0x18, 0x20, 0x58, 0x03, 0x27, 0x15,
	0x18, 0x00, 0x28, 0x25, 0x22, 0x08, 0x2D, 0x21, 0x28, 0x19, 0x2C, 0x12,
	0x15, 0x1A, 0x0B, 0x5A, 0x58, 0x76, 0x22, 0x36, 0x1E, 0x1C, 0x14, 0x3F,
	0x18, 0x0D, 0x1C, 0x29, 0x0A, 0x2C, 0x24, 0x09, 0x6D, 0x3A, 0x03, 0x3E,
	0x29, 0x69, 0x3E, 0x18, 0x3F, 0x1D, 0x23, 0x20, 0x52, 0x0A, 0x13, 0x34,
	0x2E, 0x2B, 0x03, 0x2C, 0x13, 0x25, 0x2D, 0x2C, 0x04, 0x04, 0x01, 0x12,
	0x38, 0x5B, 0x32, 0x3F, 0x3B, 0x06, 0x1D, 0x08, 0x24, 0x23, 0x2D, 0x0A,
	0x77, 0x2F, 0x00, 0x5A, 0x11, 0x2B, 0x5E, 0x24, 0x5D, 0x28, 0x37, 0x5C,
	0x57, 0x21, 0x59, 0x07, 0x1E, 0x23, 0x3A, 0x18, 0x7B, 0x5B, 0x16, 0x5F,
	0x3B, 0x24, 0x00, 0x33, 0x27, 0x5B, 0x24, 0x04, 0x2E, 0x09, 0x53, 0x11,
	0x21, 0x0A, 0x41, 0x32, 0x07, 0x03, 0x59, 0x3F, 0x53, 0x29, 0x0B, 0x32,
	0x3E, 0x0E, 0x25, 0x16, 0x08, 0x19, 0x3C, 0x0A, 0x14, 0x2D, 0x06, 0x5F,
	0x6D, 0x22, 0x4E, 0x5A, 0x5A, 0x71, 0x07, 0x26, 0x27, 0x28, 0x7A, 0x2F,
	0x11, 0x27, 0x1E, 0x13, 0x5F, 0x36, 0x24, 0x5B, 0x0E, 0x1B, 0x26, 0x34,
	0x2A, 0x08, 0x2E, 0x23, 0x3F, 0x2C, 0x76, 0x3D, 0x08, 0x2B, 0x58, 0x70,
	0x01, 0x32, 0x28, 0x18, 0x25, 0x26, 0x14, 0x09, 0x5A, 0x23, 0x5E, 0x20,
	0x08, 0x29, 0x33, 0x3D, 0x2F, 0x5E, 0x3B, 0x12, 0x1A, 0x2B, 0x0A, 0x00,
	0x7B, 0x03, 0x09, 0x27, 0x5D, 0x13, 0x47, 0x06, 0x5F, 0x33, 0x7A, 0x28,
	0x59, 0x00, 0x1F, 0x01, 0x18, 0x0E, 0x00, 0x32, 0x38, 0x1D, 0x33, 0x1A,
	0x1D, 0x31, 0x14, 0x22, 0x3F, 0x20, 0x76, 0x2A, 0x3B, 0x2F, 0x28, 0x13,
	0x5B, 0x38, 0x3F, 0x18, 0x04, 0x16, 0x52, 0x56, 0x2E, 0x3B, 0x2E, 0x1B,
	0x03, 0x21, 0x00, 0x59, 0x30, 0x1D, 0x52, 0x6D, 0x36, 0x54, 0x1B, 0x1E,
	0x2F, 0x09, 0x13, 0x5E, 0x0E, 0x15, 0x0B, 0x50, 0x57, 0x06, 0x7B, 0x59,
	0x35, 0x0D, 0x58, 0x05, 0x39, 0x17, 0x1C, 0x02, 0x31, 0x21, 0x10, 0x2C,
	0x19, 0x36, 0x3C, 0x08, 0x1B, 0x11, 0x6D, 0x1E, 0x03, 0x41, 0x5A, 0x15,
	0x05, 0x16, 0x28, 0x31, 0x06, 0x0F, 0x09, 0x58, 0x3A, 0x0E, 0x35, 0x35,
	0x1D, 0x07, 0x75, 0x0F, 0x55, 0x3A, 0x12, 0x1B, 0x55, 0x39, 0x34, 0x29,
	0x33, 0x5F, 0x59, 0x2F, 0x5E, 0x06, 0x1F, 0x22, 0x5A, 0x39, 0x2A, 0x25,
	0x25, 0x0F, 0x11, 0x09, 0x04, 0x57, 0x26, 0x3D, 0x10, 0x08, 0x07, 0x59,
	0x12, 0x0A, 0x23, 0x14, 0x3A, 0x53, 0x69, 0x20, 0x50, 0x23, 0x03, 0x17,
	0x07, 0x2E, 0x05, 0x28, 0x77, 0x2F, 0x11, 0x2F, 0x1A, 0x2D, 0x2E, 0x02,
	0x2A, 0x53, 0x2A, 0x24, 0x20, 0x08, 0x00, 0x2B, 0x25, 0x28, 0x0D, 0x21,
	0x0D, 0x3F, 0x22, 0x45, 0x53, 0x2C, 0x29, 0x09, 0x5E, 0x5A, 0x27, 0x1D,
	0x2F, 0x04, 0x01, 0x15, 0x1F, 0x51, 0x0A, 0x53, 0x2C, 0x36, 0x4E, 0x2F,
	0x0F, 0x1A, 0x58, 0x29, 0x17, 0x24, 0x0C, 0x19, 0x59, 0x24, 0x2D, 0x08,
	0x0B, 0x27, 0x16, 0x5D, 0x25, 0x5A, 0x57, 0x28, 0x00, 0x34, 0x0E, 0x54,
	0x0F, 0x5B, 0x05, 0x01, 0x04, 0x01, 0x24, 0x24, 0x20, 0x03, 0x34, 0x2D,
	0x3B, 0x27, 0x08, 0x0D, 0x05, 0x07, 0x1E, 0x05, 0x1F, 0x12, 0x74, 0x58,
	0x24, 0x58, 0x5E, 0x38, 0x2E, 0x18, 0x2F, 0x3B, 0x03, 0x3C, 0x28, 0x04,
	0x3A, 0x31, 0x0D, 0x2D, 0x5F, 0x0D, 0x6D, 0x24, 0x03, 0x41, 0x0F, 0x2E,
	0x02, 0x06, 0x08, 0x22, 0x3B, 0x1B, 0x23, 0x34, 0x28, 0x17, 0x0B, 0x2B,
	0x05, 0x24, 0x20, 0x5E, 0x58, 0x21, 0x3A, 0x10, 0x03, 0x55, 0x5F, 0x29,
	0x77, 0x00, 0x53, 0x2F, 0x44, 0x06, 0x5C, 0x09, 0x58, 0x5F, 0x15, 0x2A,
	0x4E, 0x5A, 0x53, 0x25, 0x0F, 0x53, 0x16, 0x5C, 0x27, 0x01, 0x00, 0x34,
	0x39, 0x34, 0x59, 0x1B, 0x0B, 0x58, 0x30, 0x47, 0x14, 0x5E, 0x09, 0x0D,
	0x3D, 0x10, 0x1D, 0x05, 0x34, 0x54, 0x50, 0x26, 0x33, 0x25, 0x38, 0x28,
	0x25, 0x1C, 0x05, 0x59, 0x0C, 0x1E, 0x2F, 0x0C, 0x25, 0x09, 0x1B, 0x11,
	0x7A, 0x0E, 0x03, 0x5E, 0x52, 0x05, 0x09, 0x2F, 0x0C, 0x22, 0x14, 0x3B,
	0x56, 0x19, 0x23, 0x29, 0x0F, 0x55, 0x2F, 0x08, 0x00, 0x23, 0x35, 0x1C,
	0x0C, 0x12, 0x15, 0x34, 0x05, 0x20, 0x72, 0x05, 0x51, 0x18, 0x3E, 0x13,
	0x15, 0x31, 0x16, 0x39, 0x0B, 0x27, 0x0E, 0x3D, 0x28, 0x73, 0x01, 0x2C,
	0x18, 0x2D, 0x07, 0x5C, 0x0B, 0x0B, 0x3E, 0x69, 0x54, 0x4A, 0x5F, 0x40,
	0x33, 0x55, 0x0D, 0x18, 0x07, 0x74, 0x5F, 0x22, 0x0B, 0x1F, 0x2E, 0x07,
	0x23, 0x3C, 0x0E, 0x11, 0x3A, 0x0B, 0x5E, 0x00, 0x72, 0x15, 0x31, 0x37,
	0x22, 0x75, 0x06, 0x2E, 0x5C, 0x1C, 0x2B, 0x26, 0x09, 0x36, 0x58, 0x76,
	0x27, 0x34, 0x25, 0x5D, 0x3A, 0x3B, 0x08, 0x58, 0x2C, 0x73, 0x1E, 0x58,
	0x0D, 0x38, 0x3B, 0x54, 0x25, 0x34, 0x29, 0x77, 0x2D, 0x2B, 0x2A, 0x1D,
	0x03, 0x3C, 0x28, 0x14, 0x3A, 0x01, 0x59, 0x55, 0x06, 0x5F, 0x7B, 0x21,
	0x20, 0x45, 0x3A, 0x3B, 0x3D, 0x23, 0x37, 0x2F, 0x21, 0x06, 0x34, 0x09,
	0x2A, 0x76, 0x2F, 0x59, 0x29, 0x5E, 0x03, 0x3C, 0x20, 0x5D, 0x22, 0x20,
	0x25, 0x2B, 0x56, 0x29, 0x77, 0x26, 0x59, 0x2B, 0x1C, 0x30, 0x02, 0x2F,
	0x0F, 0x2F, 0x14, 0x55, 0x23, 0x5F, 0x1A, 0x26, 0x2E, 0x14, 0x3F, 0x08,
	0x0B, 0x39, 0x51, 0x16, 0x2D, 0x38, 0x16, 0x14, 0x3C, 0x07, 0x6D, 0x01,
	0x36, 0x37, 0x28, 0x7A, 0x2E, 0x2B, 0x2D, 0x31, 0x25, 0x20, 0x16, 0x21,
	0x00, 0x09, 0x1F, 0x23, 0x58, 0x38, 0x26, 0x07, 0x0F, 0x5F, 0x0C, 0x30,
	0x2B, 0x30, 0x3D, 0x31, 0x05, 0x1B, 0x29, 0x5B, 0x02, 0x07, 0x28, 0x28,
	0x07, 0x01, 0x0C, 0x1E, 0x38, 0x1F, 0x5C, 0x0F, 0x3C, 0x32, 0x3C, 0x11,
	0x11, 0x22, 0x3B, 0x08, 0x03, 0x27, 0x18, 0x59, 0x45, 0x53, 0x20, 0x5C,
	0x15, 0x28, 0x1C, 0x14, 0x25, 0x51, 0x1F, 0x59, 0x29, 0x0D, 0x30, 0x17,
	0x21, 0x74, 0x24, 0x37, 0x0C, 0x1C, 0x25, 0x59, 0x2B, 0x1B, 0x5C, 0x77,
	0x1B, 0x0F, 0x08, 0x5D, 0x14, 0x34, 0x03, 0x41, 0x2D, 0x27, 0x0E, 0x35,
	0x56, 0x0E, 0x6D, 0x5C, 0x0A, 0x0F, 0x06, 0x03, 0x20, 0x20, 0x39, 0x00,
	0x00, 0x21, 0x06, 0x03, 0x3A, 0x05, 0x58, 0x30, 0x3D, 0x2F, 0x37, 0x16,
	0x27, 0x1D, 0x04, 0x37, 0x0D, 0x29, 0x3B, 0x2A, 0x29, 0x2B, 0x59, 0x2D,
	0x08, 0x2A, 0x15, 0x30, 0x36, 0x1C, 0x0E, 0x15, 0x3B, 0x5E, 0x28, 0x27,
	0x47, 0x10, 0x59, 0x5B, 0x16, 0x2A, 0x2A, 0x20, 0x1D, 0x12, 0x2E, 0x05,
	0x18, 0x18, 0x3A, 0x2F, 0x30, 0x05, 0x5F, 0x09, 0x47, 0x56, 0x05, 0x2E,
	0x0F, 0x06, 0x37, 0x2F, 0x44, 0x25, 0x0D, 0x30, 0x26, 0x3A, 0x0E, 0x04,
	0x39, 0x34, 0x2A, 0x76, 0x2F, 0x0C, 0x5A, 0x05, 0x2F, 0x34, 0x0A, 0x36,
	0x1E, 0x36, 0x1E, 0x55, 0x01, 0x2C, 0x2B, 0x00, 0x37, 0x18, 0x0A, 0x0E,
	0x43, 0x0E, 0x1C, 0x11, 0x73, 0x58, 0x29, 0x1C, 0x03, 0x76, 0x3F, 0x2C,
	0x2B, 0x0F, 0x6D, 0x55, 0x17, 0x5E, 0x2F, 0x2F, 0x18, 0x55, 0x2F, 0x53,
	0x7A, 0x08, 0x53, 0x2D, 0x38, 0x69, 0x5E, 0x33, 0x2A, 0x1C, 0x34, 0x22,
	0x3B, 0x22, 0x0A, 0x33, 0x2A, 0x3B, 0x1B, 0x29, 0x30, 0x02, 0x1B, 0x09,
	0x1F, 0x32, 0x1C, 0x20, 0x1C, 0x08, 0x76, 0x26, 0x4E, 0x5D, 0x3F, 0x33,
	0x19, 0x4E, 0x5E, 0x19, 0x38, 0x1B, 0x29, 0x05, 0x1F, 0x1B, 0x2E, 0x02,
	0x3C, 0x53, 0x2A, 0x28, 0x16, 0x07, 0x1E, 0x32, 0x29, 0x2D, 0x24, 0x3D,
	0x74, 0x22, 0x55, 0x5C, 0x22, 0x11, 0x0F, 0x2D, 0x37, 0x18, 0x72, 0x23,
	0x13, 0x18, 0x25, 0x08, 0x3D, 0x0E, 0x5A, 0x06, 0x7A, 0x59, 0x04, 0x1F,
	0x03, 0x70, 0x55, 0x18, 0x28, 0x25, 0x0F, 0x5F, 0x58, 0x03, 0x3D, 0x2D,
	0x08, 0x38, 0x17, 0x3A, 0x10, 0x0E, 0x2A, 0x25, 0x25, 0x21, 0x04, 0x02,
	0x1D, 0x22, 0x12, 0x5C, 0x0B, 0x5B, 0x0C, 0x18, 0x26, 0x4A, 0x14, 0x1C,
	0x18, 0x0A, 0x55, 0x0F, 0x00, 0x09, 0x3B, 0x20, 0x1C, 0x2D, 0x1A, 0x25,
	0x04, 0x3E, 0x1E, 0x27, 0x04, 0x55, 0x1F, 0x07, 0x17, 0x04, 0x09, 0x28,
	0x00, 0x7A, 0x3B, 0x02, 0x1D, 0x0C, 0x2E, 0x0D, 0x52, 0x0C, 0x2F, 0x06,
	0x5F, 0x4E, 0x36, 0x11, 0x13, 0x39, 0x2A, 0x21, 0x02, 0x1A, 0x19, 0x4A,
	0x00, 0x31, 0x06, 0x5D, 0x55, 0x09, 0x5C, 0x34, 0x59, 0x04, 0x1D, 0x22,
	0x01, 0x47, 0x51, 0x26, 0x08, 0x0D, 0x3B, 0x29, 0x2F, 0x09, 0x2C, 0x0B,
	0x31, 0x3A, 0x5E, 0x3B, 0x29, 0x32, 0x2F, 0x1D, 0x03, 0x23, 0x30, 0x38,
	0x0C, 0x01, 0x14, 0x55, 0x04, 0x44, 0x75, 0x26, 0x12, 0x0F, 0x1C, 0x0B,
	0x3B, 0x32, 0x08, 0x1E, 0x37, 0x3D, 0x57, 0x1A, 0x44, 0x25, 0x0D, 0x30,
	0x2A, 0x1C, 0x12, 0x15, 0x04, 0x3B, 0x2F, 0x37, 0x2D, 0x4A, 0x3A, 0x23,
	0x25, 0x3C, 0x19, 0x39, 0x22, 0x07, 0x29, 0x07, 0x34, 0x53, 0x75, 0x3E,
	0x0D, 0x16, 0x29, 0x30, 0x14, 0x51, 0x45, 0x5F, 0x3B, 0x3B, 0x59, 0x5F,
	0x2E, 0x18, 0x2D, 0x39, 0x2F, 0x3B, 0x08, 0x27, 0x30, 0x27, 0x1A, 0x07,
	0x5B, 0x23, 0x0F, 0x52, 0x0C, 0x1B, 0x2A, 0x34, 0x01, 0x35, 0x2A, 0x18,
	0x24, 0x12, 0x04, 0x16, 0x19, 0x08, 0x1E, 0x77, 0x28, 0x53, 0x3D, 0x24,
	0x03, 0x0A, 0x2D, 0x22, 0x06, 0x7B, 0x26, 0x1B, 0x34, 0x01, 0x14, 0x3F,
	0x04, 0x25, 0x53, 0x34, 0x21, 0x19, 0x58, 0x3A, 0x3B, 0x35, 0x23, 0x5E,
	0x2E, 0x16, 0x26, 0x33, 0x39, 0x20, 0x21, 0x1A, 0x09, 0x5E, 0x1A, 0x7A,
	0x2F, 0x51, 0x00, 0x06, 0x0B, 0x0E, 0x0D, 0x14, 0x05, 0x08, 0x2F, 0x18,
	0x1B, 0x24, 0x21, 0x3D, 0x13, 0x18, 0x1C, 0x27, 0x3D, 0x11, 0x01, 0x02,
	0x17, 0x1A, 0x0E, 0x16, 0x3A, 0x2E, 0x0E, 0x2A, 0x0A, 0x33, 0x0C, 0x2F,
	0x0B, 0x01, 0x00, 0x71, 0x08, 0x11, 0x2D, 0x3A, 0x32, 0x39, 0x28, 0x00,
	0x0D, 0x00, 0x19, 0x14, 0x18, 0x29, 0x30, 0x01, 0x13, 0x5F, 0x26, 0x25,
	0x54, 0x18, 0x0A, 0x2A, 0x2C, 0x1E, 0x31, 0x3A, 0x39, 0x70, 0x0E, 0x17,
	0x5F, 0x26, 0x38, 0x1C, 0x4A, 0x28, 0x1B, 0x07, 0x15, 0x22, 0x3A, 0x13,
	0x1A, 0x2B, 0x14, 0x09, 0x5A, 0x10, 0x2D, 0x09, 0x2C, 0x13, 0x09, 0x36,
	0x37, 0x1E, 0x23, 0x0C, 0x16, 0x29, 0x0F, 0x58, 0x2E, 0x24, 0x0C, 0x00,
	0x0A, 0x04, 0x39, 0x00, 0x25, 0x27, 0x18, 0x1B, 0x0F, 0x45, 0x53, 0x36,
	0x0F, 0x2E, 0x39, 0x5C, 0x01, 0x20, 0x0D, 0x36, 0x01, 0x0D, 0x34, 0x56,
	0x3F, 0x0E, 0x18, 0x0E, 0x09, 0x27, 0x1C, 0x10, 0x5F, 0x15, 0x57, 0x21,
	0x29, 0x3C, 0x0A, 0x57, 0x22, 0x07, 0x55, 0x54, 0x26, 0x5C, 0x73, 0x02,
	0x51, 0x0B, 0x19, 0x77, 0x5B, 0x4E, 0x20, 0x07, 0x18, 0x04, 0x2B, 0x17,
	0x3E, 0x07, 0x3F, 0x36, 0x22, 0x0C, 0x27, 0x36, 0x0D, 0x0B, 0x52, 0x0E,
	0x38, 0x59, 0x36, 0x38, 0x11, 0x2A, 0x39, 0x27, 0x29, 0x07, 0x22, 0x02,
	0x2B, 0x3C, 0x70, 0x03, 0x31, 0x2B, 0x44, 0x37, 0x2A, 0x09, 0x3F, 0x12,
	0x08, 0x07, 0x07, 0x0F, 0x1A, 0x35, 0x00, 0x4E, 0x2D, 0x53, 0x2C, 0x1F,
	0x27, 0x5D, 0x5A, 0x31, 0x20, 0x56, 0x2C, 0x44, 0x28, 0x1C, 0x20, 0x1E,
	0x26, 0x2D, 0x26, 0x29, 0x17, 0x23, 0x20, 0x3E, 0x07, 0x5E, 0x5E, 0x03,
	0x1D, 0x56, 0x21, 0x2A, 0x1A, 0x3C, 0x33, 0x45, 0x06, 0x32, 0x1A, 0x27,
	0x0A, 0x3D, 0x75, 0x54, 0x07, 0x02, 0x52, 0x2F, 0x20, 0x08, 0x2C, 0x19,
	0x03, 0x27, 0x0A, 0x3C, 0x08, 0x2B, 0x28, 0x2F, 0x21, 0x53, 0x70, 0x21,
	0x18, 0x1A, 0x5F, 0x0D, 0x08, 0x05, 0x39, 0x1E, 0x2A, 0x47, 0x17, 0x1D,
	0x2A, 0x37, 0x3D, 0x1B, 0x09, 0x3B, 0x35, 0x16, 0x28, 0x25, 0x08, 0x03,
	0x47, 0x35, 0x5E, 0x0C, 0x29, 0x16, 0x56, 0x09, 0x22, 0x73, 0x21, 0x23,
	0x1B, 0x32, 0x3B, 0x3D, 0x16, 0x5A, 0x06, 0x73, 0x03, 0x56, 0x17, 0x1F,
	0x07, 0x1A, 0x0A, 0x59, 0x29, 0x1A, 0x08, 0x02, 0x36, 0x2A, 0x37, 0x18,
	0x10, 0x01, 0x2A, 0x0F, 0x29, 0x0F, 0x24, 0x2E, 0x27, 0x3C, 0x51, 0x08,
	0x2A, 0x32, 0x00, 0x31, 0x2D, 0x28, 0x13, 0x35, 0x08, 0x01, 0x0A, 0x28,
	0x23, 0x2A, 0x19, 0x5A, 0x10, 0x3B, 0x4A, 0x5B, 0x2D, 0x73, 0x03, 0x05,
	0x2C, 0x40, 0x13, 0x5F, 0x06, 0x2A, 0x13, 0x70, 0x00, 0x55, 0x57, 0x26,
	0x03, 0x5E, 0x30, 0x06, 0x22, 0x14, 0x23, 0x27, 0x1C, 0x0D, 0x14, 0x2B,
	0x0A, 0x25, 0x05, 0x36, 0x5C, 0x08, 0x08, 0x1B, 0x32, 0x2E, 0x39, 0x41,
	0x1F, 0x2D, 0x28, 0x2C, 0x2A, 0x00, 0x0E, 0x5E, 0x08, 0x34, 0x2D, 0x3B,
	0x21, 0x18, 0x28, 0x5C, 0x3A, 0x2A, 0x13, 0x5C, 0x31, 0x74, 0x28, 0x37,
	0x37, 0x3E, 0x01, 0x47, 0x35, 0x56, 0x0C, 0x2A, 0x35, 0x36, 0x08, 0x40,
	0x01, 0x01, 0x30, 0x0B, 0x52, 0x7A, 0x24, 0x51, 0x5D, 0x2E, 0x2F, 0x22,
	0x31, 0x27, 0x24, 0x13, 0x23, 0x55, 0x3D, 0x3C, 0x37, 0x3C, 0x08, 0x2A,
	0x0D, 0x33, 0x18, 0x27, 0x09, 0x29, 0x13, 0x2E, 0x08, 0x3F, 0x2D, 0x77,
	0x23, 0x18, 0x2B, 0x23, 0x3A, 0x3B, 0x08, 0x58, 0x29, 0x15, 0x3D, 0x4A,
	0x3C, 0x53, 0x2B, 0x07, 0x19, 0x23, 0x5C, 0x29, 0x3F, 0x24, 0x5A, 0x21,
	0x0B, 0x1A, 0x4E, 0x5D, 0x3A, 0x74, 0x1A, 0x17, 0x2F, 0x44, 0x08, 0x20,
	0x30, 0x2C, 0x5C, 0x6D, 0x25, 0x03, 0x24, 0x00, 0x3A, 0x25, 0x1B, 0x5C,
	0x05, 0x03, 0x43, 0x54, 0x23, 0x02, 0x7A, 0x2B, 0x54, 0x28, 0x3C, 0x03,
	0x1E, 0x22, 0x38, 0x00, 0x28, 0x3C, 0x06, 0x58, 0x22, 0x21, 0x19, 0x28,
	0x0B, 0x3C, 0x21, 0x38, 0x28, 0x3F, 0x40, 0x0B, 0x43, 0x31, 0x02, 0x58,
	0x35, 0x34, 0x34, 0x45, 0x2A, 0x31, 0x0B, 0x58, 0x09, 0x3B, 0x35, 0x38,
	0x28, 0x2A, 0x53, 0x29, 0x59, 0x22, 0x2B, 0x39, 0x71, 0x34, 0x52, 0x56,
	0x03, 0x69, 0x29, 0x11, 0x2F, 0x27, 0x29, 0x2F, 0x0A, 0x28, 0x3C, 0x07,
	0x24, 0x23, 0x26, 0x59, 0x24, 0x26, 0x26, 0x3F, 0x20, 0x13, 0x27, 0x2B,
	0x01, 0x0F, 0x1A, 0x5B, 0x20, 0x22, 0x00, 0x26, 0x07, 0x20, 0x21, 0x2A,
	0x0A, 0x2D, 0x03, 0x05, 0x59, 0x76, 0x28, 0x59, 0x06, 0x21, 0x06, 0x38,
	0x38, 0x07, 0x44, 0x27, 0x24, 0x51, 0x2A, 0x06, 0x7A, 0x38, 0x07, 0x59,
	0x12, 0x03, 0x3E, 0x20, 0x5B, 0x0C, 0x01, 0x15, 0x0F, 0x24, 0x28, 0x3A,
	0x35, 0x12, 0x34, 0x0D, 0x13, 0x58, 0x06, 0x57, 0x5B, 0x72, 0x5C, 0x0B,
	0x2A, 0x3C, 0x28, 0x5D, 0x2F, 0x05, 0x2F, 0x70, 0x2D, 0x07, 0x25, 0x3B,
	0x25, 0x24, 0x18, 0x0C, 0x00, 0x05, 0x5D, 0x08, 0x00, 0x21, 0x76, 0x2B,
	0x0C, 0x3A, 0x53, 0x00, 0x54, 0x13, 0x3C, 0x09, 0x74, 0x26, 0x12, 0x25,
	0x38, 0x70, 0x0E, 0x14, 0x22, 0x09, 0x75, 0x21, 0x37, 0x37, 0x29, 0x17,
	0x2D, 0x05, 0x05, 0x2C, 0x3B, 0x29, 0x02, 0x24, 0x02, 0x1B, 0x3B, 0x58,
	0x56, 0x33, 0x2F, 0x3D, 0x4A, 0x3D, 0x04, 0x25, 0x43, 0x18, 0x0F, 0x3A,
	0x2D, 0x2E, 0x55, 0x21, 0x18, 0x14, 0x3B, 0x56, 0x36, 0x44, 0x16, 0x02,
	0x0A, 0x17, 0x39, 0x38, 0x3F, 0x2D, 0x14, 0x3D, 0x1A, 0x54, 0x23, 0x5F,
	0x13, 0x2C, 0x58, 0x24, 0x00, 0x03, 0x11, 0x3D, 0x08, 0x19, 0x2D, 0x77,
	0x26, 0x32, 0x2C, 0x1D, 0x00, 0x2F, 0x30, 0x39, 0x38, 0x08, 0x43, 0x3B,
	0x5F, 0x3B, 0x27, 0x3D, 0x53, 0x20, 0x05, 0x74, 0x3A, 0x11, 0x27, 0x31,
	0x0E, 0x5D, 0x38, 0x2A, 0x3B, 0x35, 0x34, 0x39, 0x21, 0x38, 0x11, 0x3D,
	0x30, 0x29, 0x53, 0x13, 0x27, 0x38, 0x19, 0x33, 0x7A, 0x54, 0x39, 0x5D,
	0x04, 0x26, 0x34, 0x4E, 0x2F, 0x3C, 0x16, 0x21, 0x13, 0x0A, 0x3F, 0x0E,
	0x04, 0x36, 0x34, 0x5C, 0x71, 0x1D, 0x52, 0x19, 0x33, 0x0B, 0x2F, 0x12,
	0x27, 0x1E, 0x11, 0x21, 0x51, 0x2D, 0x3F, 0x30, 0x3D, 0x00, 0x34, 0x2C,
	0x3B, 0x29, 0x10, 0x16, 0x13, 0x30, 0x1D, 0x37, 0x05, 0x29, 0x2E, 0x2F,
	0x20, 0x5D, 0x12, 0x17, 0x1E, 0x18, 0x3E, 0x32, 0x34, 0x1B, 0x25, 0x36,
	0x40, 0x13, 0x35, 0x06, 0x41, 0x1C, 0x0A, 0x25, 0x56, 0x19, 0x2D, 0x77,
	0x26, 0x09, 0x57, 0x0D, 0x09, 0x47, 0x00, 0x2D, 0x07, 0x69, 0x5F, 0x53,
	0x34, 0x3D, 0x76, 0x2A, 0x18, 0x2A, 0x3C, 0x03, 0x18, 0x20, 0x26, 0x31,
	0x03, 0x0F, 0x08, 0x1A, 0x0C, 0x0A, 0x1B, 0x00, 0x05, 0x3B, 0x31, 0x2D,
	0x4A, 0x3A, 0x2E, 0x2A, 0x5D, 0x34, 0x3C, 0x19, 0x73, 0x0E, 0x3B, 0x05,
	0x39, 0x21, 0x22, 0x4A, 0x06, 0x1F, 0x2F, 0x16, 0x02, 0x24, 0x59, 0x0E,
	0x3C, 0x14, 0x01, 0x01, 0x38, 0x15, 0x27, 0x05, 0x1B, 0x1A, 0x06, 0x31,
	0x1C, 0x1C, 0x01, 0x36, 0x37, 0x37, 0x2A, 0x07, 0x0B, 0x26, 0x19, 0x2A,
	0x77, 0x2D, 0x00, 0x2C, 0x1F, 0x0F, 0x27, 0x09, 0x2D, 0x1B, 0x69, 0x28,
	0x14, 0x28, 0x39, 0x07, 0x3C, 0x26, 0x58, 0x29, 0x14, 0x02, 0x02, 0x2A,
	0x53, 0x2D, 0x2E, 0x20, 0x45, 0x07, 0x33, 0x04, 0x36, 0x07, 0x53, 0x7B,
	0x20, 0x15, 0x0A, 0x07, 0x2D, 0x22, 0x37, 0x2A, 0x03, 0x0D, 0x1B, 0x32,
	0x21, 0x1E, 0x07, 0x3E, 0x0A, 0x26, 0x05, 0x7A, 0x14, 0x52, 0x14, 0x00,
	0x74, 0x35, 0x22, 0x56, 0x28, 0x08, 0x28, 0x54, 0x09, 0x3B, 0x13, 0x20,
	0x3B, 0x20, 0x2A, 0x15, 0x2F, 0x19, 0x37, 0x12, 0x20, 0x36, 0x00, 0x34,
	0x5E, 0x36, 0x5B, 0x1B, 0x57, 0x32, 0x13, 0x0F, 0x24, 0x18, 0x1B, 0x35,
	0x20, 0x50, 0x14, 0x5E, 0x23, 0x58, 0x20, 0x0D, 0x21, 0x70, 0x3F, 0x52,
	0x03, 0x27, 0x7B, 0x23, 0x22, 0x16, 0x06, 0x0D, 0x22, 0x05, 0x02, 0x25,
	0x0C, 0x0F, 0x54, 0x5D, 0x44, 0x75, 0x0B, 0x13, 0x1D, 0x59, 0x10, 0x04,
	0x34, 0x29, 0x53, 0x72, 0x01, 0x0B, 0x21, 0x07, 0x38, 0x20, 0x2F, 0x27,
	0x5E, 0x30, 0x06, 0x16, 0x58, 0x2C, 0x69, 0x2A, 0x07, 0x3D, 0x5F, 0x1A,
	0x0A, 0x1B, 0x19, 0x52, 0x10, 0x3A, 0x0E, 0x04, 0x07, 0x71, 0x5F, 0x02,
	0x02, 0x5A, 0x2C, 0x14, 0x02, 0x3A, 0x5E, 0x1A, 0x15, 0x05, 0x38, 0x39,
	0x20, 0x1B, 0x22, 0x34, 0x24, 0x2B, 0x2E, 0x17, 0x5B, 0x3D, 0x23, 0x2F,
	0x4E, 0x39, 0x0A, 0x13, 0x19, 0x30, 0x21, 0x3A, 0x0E, 0x1B, 0x0A, 0x05,
	0x2C, 0x0F, 0x16, 0x00, 0x3A, 0x44, 0x10, 0x3C, 0x51, 0x21, 0x04, 0x0A,
	0x0B, 0x25, 0x19, 0x26, 0x3B, 0x20, 0x31, 0x5C, 0x40, 0x0F, 0x04, 0x12,
	0x3F, 0x06, 0x76, 0x3B, 0x57, 0x57, 0x3F, 0x0E, 0x04, 0x34, 0x14, 0x08,
	0x2B, 0x25, 0x17, 0x38, 0x1C, 0x0C, 0x54, 0x23, 0x1D, 0x39, 0x23, 0x19,
	0x12, 0x5B, 0x2C, 0x13, 0x1F, 0x51, 0x27, 0x0D, 0x20, 0x05, 0x03, 0x05,
	0x39, 0x2F, 0x2B, 0x1B, 0x18, 0x39, 0x36, 0x0D, 0x31, 0x3C, 0x1D, 0x70,
	0x03, 0x58, 0x5C, 0x5D, 0x3A, 0x55, 0x4A, 0x41, 0x44, 0x00, 0x00, 0x0E,
	0x57, 0x3A, 0x03, 0x0B, 0x52, 0x19, 0x23, 0x29, 0x26, 0x55, 0x2A, 0x53,
	0x0C, 0x15, 0x22, 0x3E, 0x1E, 0x21, 0x5D, 0x29, 0x00, 0x00, 0x2C, 0x25,
	0x05, 0x1B, 0x23, 0x7B, 0x1A, 0x34, 0x22, 0x22, 0x74, 0x2E, 0x2C, 0x1E,
	0x5D, 0x0B, 0x5E, 0x2B, 0x5C, 0x0E, 0x30, 0x3A, 0x02, 0x24, 0x5B, 0x03,
	0x07, 0x24, 0x28, 0x2A, 0x36, 0x0B, 0x2F, 0x17, 0x20, 0x24, 0x38, 0x2C,
	0x3A, 0x5F, 0x0E, 0x21, 0x28, 0x3B, 0x27, 0x70, 0x05, 0x2B, 0x00, 0x13,
	0x32, 0x15, 0x25, 0x14, 0x53, 0x05, 0x5F, 0x11, 0x39, 0x08, 0x6D, 0x2B,
	0x50, 0x18, 0x04, 0x07, 0x43, 0x34, 0x41, 0x26, 0x0F, 0x00, 0x2C, 0x41,
	0x5F, 0x20, 0x08, 0x00, 0x2C, 0x2E, 0x25, 0x3E, 0x0A, 0x2C, 0x18, 0x00,
	0x47, 0x30, 0x3F, 0x0C, 0x1A, 0x1B, 0x35, 0x05, 0x0A, 0x77, 0x43, 0x30,
	0x3E, 0x11, 0x2F, 0x0D, 0x0F, 0x5B, 0x29, 0x08, 0x0F, 0x0E, 0x0D, 0x5A,
	0x36, 0x2E, 0x11, 0x14, 0x1E, 0x76, 0x43, 0x59, 0x20, 0x38, 0x03, 0x1A,
	0x20, 0x45, 0x39, 0x11, 0x0B, 0x34, 0x3C, 0x03, 0x71, 0x22, 0x17, 0x1B,
	0x04, 0x7B, 0x29, 0x15, 0x57, 0x3B, 0x0C, 0x3F, 0x00, 0x3E, 0x3E, 0x2F,
	0x3D, 0x2F, 0x1F, 0x2E, 0x2C, 0x2E, 0x33, 0x58, 0x5C, 0x0D, 0x21, 0x06,
	0x56, 0x5B, 0x14, 0x2D, 0x17, 0x05, 0x23, 0x0B, 0x2D, 0x00, 0x26, 0x23,
	0x34, 0x0B, 0x02, 0x17, 0x1D, 0x35, 0x36, 0x0A, 0x19, 0x07, 0x76, 0x0A,
	0x04, 0x3C, 0x5F, 0x25, 0x5C, 0x16, 0x2A, 0x1B, 0x00, 0x19, 0x33, 0x5F,
	0x0C, 0x12, 0x3D, 0x33, 0x23, 0x00, 0x14, 0x54, 0x58, 0x59, 0x0E, 0x06,
	0x16, 0x2F, 0x56, 0x29, 0x21, 0x04, 0x59, 0x09, 0x58, 0x35, 0x20, 0x0A,
	0x3E, 0x1C, 0x07, 0x59, 0x22, 0x56, 0x01, 0x20, 0x35, 0x2E, 0x5B, 0x40,
	0x7A, 0x18, 0x4E, 0x5B, 0x12, 0x12, 0x21, 0x2B, 0x39, 0x38, 0x75, 0x09,
	0x53, 0x2C, 0x12, 0x13, 0x19, 0x30, 0x58, 0x3A, 0x06, 0x35, 0x20, 0x23,
	0x2A, 0x2C, 0x27, 0x35, 0x3F, 0x25, 0x2B, 0x5E, 0x10, 0x2A, 0x08, 0x09,
	0x04, 0x30, 0x2B, 0x39, 0x38, 0x5B, 0x16, 0x0A, 0x3C, 0x2C, 0x5C, 0x04,
	0x05, 0x28, 0x0F, 0x2F, 0x2A, 0x0D, 0x32, 0x0C, 0x18, 0x3B, 0x1A, 0x13,
	0x2F, 0x59, 0x08, 0x1E, 0x3F, 0x72, 0x2F, 0x13, 0x23, 0x5F, 0x00, 0x0F,
	0x4A, 0x2B, 0x00, 0x24, 0x09, 0x35, 0x01, 0x0C, 0x29, 0x1B, 0x26, 0x34,
	0x29, 0x31, 0x05, 0x13, 0x2D, 0x20, 0x29, 0x27, 0x29, 0x08, 0x3E, 0x05,
	0x07, 0x23, 0x00, 0x5F, 0x32, 0x3C, 0x57, 0x04, 0x5A, 0x37, 0x1D, 0x37,
	0x14, 0x2F, 0x1A, 0x3B, 0x57, 0x58, 0x23, 0x14, 0x20, 0x38, 0x3C, 0x26,
	0x07, 0x2A, 0x07, 0x0B, 0x2F, 0x38, 0x26, 0x17, 0x29, 0x40, 0x0F, 0x06,
	0x58, 0x5A, 0x3B, 0x0F, 0x28, 0x16, 0x2F, 0x5E, 0x00, 0x0F, 0x0B, 0x18,
	0x53, 0x0C, 0x07, 0x4E, 0x2C, 0x08, 0x7B, 0x23, 0x18, 0x2D, 0x07, 0x2A,
	0x5B, 0x03, 0x16, 0x38, 0x3B, 0x20, 0x23, 0x38, 0x18, 0x06, 0x29, 0x02,
	0x04, 0x06, 0x11, 0x1E, 0x50, 0x56, 0x21, 0x73, 0x25, 0x0A, 0x2D, 0x59,
	0x07, 0x55, 0x28, 0x3B, 0x0E, 0x13, 0x5B, 0x17, 0x2F, 0x5E, 0x2F, 0x55,
	0x06, 0x20, 0x1C, 0x06, 0x15, 0x25, 0x56, 0x2F, 0x21, 0x03, 0x10, 0x3F,
	0x0D, 0x27, 0x27, 0x04, 0x41, 0x1C, 0x13, 0x15, 0x1B, 0x59, 0x01, 0x06,
	0x3E, 0x57, 0x37, 0x28, 0x0F, 0x1C, 0x04, 0x3F, 0x2A, 0x14, 0x07, 0x07,
	0x2F, 0x2C, 0x10, 0x2F, 0x30, 0x03, 0x5F, 0x15, 0x43, 0x35, 0x05, 0x06,
	0x18, 0x26, 0x13, 0x3F, 0x1A, 0x7B, 0x19, 0x06, 0x5F, 0x0D, 0x31, 0x26,
	0x0C, 0x3D, 0x2E, 0x72, 0x5E, 0x53, 0x5C, 0x2E, 0x71, 0x2F, 0x27, 0x5C,
	0x5A, 0x26, 0x5D, 0x25, 0x17, 0x2C, 0x13, 0x14, 0x05, 0x5D, 0x53, 0x26,
	0x1E, 0x17, 0x20, 0x19, 0x13, 0x2F, 0x56, 0x5A, 0x1F, 0x0B, 0x55, 0x2C,
	0x2F, 0x2C, 0x13, 0x27, 0x28, 0x3E, 0x26, 0x08, 0x01, 0x32, 0x0B, 0x53,
	0x72, 0x0E, 0x37, 0x2D, 0x21, 0x2D, 0x1C, 0x03, 0x58, 0x06, 0x3B, 0x01,
	0x20, 0x34, 0x2C, 0x2C, 0x2A, 0x59, 0x20, 0x5A, 0x71, 0x07, 0x31, 0x27,
	0x3D, 0x05, 0x24, 0x27, 0x08, 0x3A, 0x10, 0x07, 0x56, 0x09, 0x09, 0x29,
	0x5E, 0x55, 0x2F, 0x53, 0x01, 0x21, 0x0B, 0x18, 0x28, 0x1A, 0x00, 0x24,
	0x04, 0x22, 0x36, 0x14, 0x05, 0x5B, 0x20, 0x14, 0x07, 0x13, 0x16, 0x2F,
	0x15, 0x14, 0x07, 0x06, 0x1E, 0x12, 0x0B, 0x36, 0x08, 0x5B, 0x17, 0x15,
	0x00, 0x56, 0x3D, 0x38, 0x1A, 0x38, 0x3D, 0x3A, 0x2E, 0x0E, 0x28, 0x21,
	0x11, 0x08, 0x5C, 0x4A, 0x5F, 0x59, 0x31, 0x26, 0x0C, 0x3D, 0x12, 0x2B,
	0x29, 0x20, 0x5C, 0x3A, 0x70, 0x3D, 0x29, 0x27, 0x09, 0x1B, 0x3D, 0x02,
	0x3D, 0x1A, 0x76, 0x54, 0x00, 0x28, 0x40, 0x18, 0x07, 0x31, 0x05, 0x26,
	0x36, 0x20, 0x10, 0x08, 0x00, 0x04, 0x06, 0x51, 0x02, 0x05, 0x7A, 0x3E,
	0x2C, 0x06, 0x11, 0x00, 0x5A, 0x53, 0x1B, 0x5B, 0x34, 0x2A, 0x18, 0x1D,
	0x33, 0x7A, 0x26, 0x50, 0x16, 0x1F, 0x75, 0x00, 0x28, 0x1E, 0x11, 0x14,
	0x1F, 0x23, 0x03, 0x12, 0x07, 0x3A, 0x54, 0x25, 0x26, 0x34, 0x3C, 0x24,
	0x1D, 0x53, 0x69, 0x55, 0x18, 0x59, 0x44, 0x0D, 0x2F, 0x0A, 0x2A, 0x0E,
	0x0B, 0x2E, 0x23, 0x04, 0x5F, 0x21, 0x47, 0x33, 0x23, 0x01, 0x14, 0x03,
	0x58, 0x38, 0x31, 0x03, 0x5F, 0x06, 0x36, 0x22, 0x18, 0x1B, 0x29, 0x5B,
	0x26, 0x2B, 0x29, 0x35, 0x3C, 0x0D, 0x6D, 0x59, 0x2F, 0x1D, 0x01, 0x7A,
	0x02, 0x2B, 0x2C, 0x5C, 0x3A, 0x38, 0x02, 0x0A, 0x18, 0x7A, 0x47, 0x39,
	0x03, 0x3A, 0x16, 0x25, 0x2F, 0x2B, 0x2A, 0x37, 0x2E, 0x4A, 0x3F, 0x5D,
	0x13, 0x3C, 0x0E, 0x24, 0x06, 0x11, 0x2A, 0x57, 0x5F, 0x28, 0x23, 0x3D,
	0x14, 0x3F, 0x2C, 0x13, 0x06, 0x16, 0x2D, 0x12, 0x06, 0x59, 0x25, 0x59,
	0x28, 0x26, 0x07, 0x15, 0x0A, 0x25, 0x13, 0x26, 0x30, 0x07, 0x0A, 0x09,
	0x1E, 0x4E, 0x21, 0x44, 0x7B, 0x43, 0x0D, 0x5C, 0x40, 0x08, 0x21, 0x4A,
	0x3F, 0x44, 0x74, 0x02, 0x36, 0x2A, 0x1E, 0x27, 0x47, 0x09, 0x00, 0x44,
	0x3B, 0x1D, 0x59, 0x2C, 0x31, 0x01, 0x5C, 0x0B, 0x19, 0x03, 0x0D, 0x43,
	0x0A, 0x34, 0x2F, 0x7B, 0x1B, 0x14, 0x21, 0x5F, 0x2C, 0x36, 0x23, 0x1E,
	0x1C, 0x29, 0x1D, 0x54, 0x2C, 0x5D, 0x75, 0x16, 0x37, 0x3B, 0x20, 0x70,
	0x2F, 0x38, 0x5D, 0x52, 0x24, 0x36, 0x20, 0x5B, 0x2A, 0x7A, 0x0B, 0x54,
	0x3F, 0x0C, 0x18, 0x29, 0x05, 0x3E, 0x08, 0x08, 0x02, 0x4E, 0x38, 0x07,
	0x08, 0x0B, 0x25, 0x17, 0x32, 0x29, 0x2D, 0x36, 0x2F, 0x58, 0x0B, 0x18,
	0x28, 0x08, 0x24, 0x07, 0x0A, 0x14, 0x5A, 0x05, 0x18, 0x25, 0x0E, 0x37,
	0x3F, 0x18, 0x2A, 0x0E, 0x1E, 0x0F, 0x23, 0x43, 0x16, 0x18, 0x19, 0x25,
	0x39, 0x0C, 0x2B, 0x5E, 0x75, 0x25, 0x30, 0x1C, 0x0D, 0x76, 0x15, 0x30,
	0x1D, 0x19, 0x01, 0x25, 0x58, 0x01, 0x23, 0x0F, 0x0A, 0x30, 0x27, 0x31,
	0x36, 0x2D, 0x04, 0x21, 0x28, 0x32, 0x00, 0x17, 0x3F, 0x0A, 0x31, 0x1E,
	0x28, 0x3B, 0x1D, 0x77, 0x3E, 0x18, 0x3D, 0x11, 0x16, 0x09, 0x30, 0x0F,
	0x44, 0x10, 0x00, 0x00, 0x3E, 0x0D, 0x14, 0x16, 0x50, 0x2C, 0x26, 0x11,
	0x06, 0x59, 0x23, 0x1B, 0x16, 0x47, 0x17, 0x27, 0x11, 0x01, 0x27, 0x3B,
	0x07, 0x0E, 0x08, 0x18, 0x39, 0x3E, 0x5F, 0x77, 0x43, 0x1B, 0x1C, 0x27,
	0x03, 0x20, 0x0D, 0x21, 0x22, 0x0A, 0x1B, 0x10, 0x2C, 0x20, 0x74, 0x3E,
	0x25, 0x3B, 0x20, 0x30, 0x2B, 0x16, 0x05, 0x5E, 0x09, 0x24, 0x13, 0x18,
	0x19, 0x11, 0x2E, 0x1B, 0x22, 0x12, 0x07, 0x3C, 0x22, 0x3D, 0x44, 0x32,
	0x3E, 0x18, 0x2A, 0x11, 0x10, 0x5C, 0x2A, 0x03, 0x28, 0x23, 0x5F, 0x4A,
	0x57, 0x3B, 0x70, 0x47, 0x1B, 0x2B, 0x18, 0x07, 0x35, 0x12, 0x58, 0x1F,
	0x7A, 0x24, 0x00, 0x39, 0x11, 0x1B, 0x2A, 0x36, 0x57, 0x53, 0x05, 0x5A,
	0x52, 0x03, 0x20, 0x13, 0x3B, 0x30, 0x00, 0x22, 0x00, 0x07, 0x25, 0x0B,
	0x3F, 0x0F, 0x0B, 0x3B, 0x56, 0x0A, 0x16, 0x1A, 0x2B, 0x1B, 0x38, 0x03,
	0x54, 0x2E, 0x16, 0x1E, 0x25, 0x5D, 0x03, 0x5D, 0x2A, 0x0A, 0x27, 0x28,
	0x05, 0x2E, 0x2C, 0x05, 0x32, 0x0C, 0x52, 0x30, 0x36, 0x29, 0x3F, 0x5A,
	0x08, 0x23, 0x55, 0x39, 0x2D, 0x3A, 0x38, 0x59, 0x08, 0x44, 0x7B, 0x2A,
	0x2C, 0x04, 0x1D, 0x04, 0x38, 0x25, 0x3A, 0x06, 0x20, 0x1E, 0x2D, 0x17,
	0x03, 0x13, 0x0E, 0x55, 0x25, 0x5B, 0x0E, 0x01, 0x22, 0x38, 0x1D, 0x2B,
	0x36, 0x39, 0x08, 0x5C, 0x75, 0x22, 0x53, 0x2F, 0x19, 0x01, 0x24, 0x0A,
	0x1B, 0x29, 0x2B, 0x3A, 0x35, 0x3B, 0x22, 0x0D, 0x05, 0x04, 0x41, 0x5A,
	0x29, 0x0E, 0x17, 0x57, 0x44, 0x08, 0x35, 0x56, 0x5A, 0x3F, 0x32, 0x0A,
	0x14, 0x38, 0x1F, 0x1A, 0x20, 0x05, 0x26, 0x3B, 0x18, 0x3A, 0x2A, 0x0C,
	0x28, 0x7B, 0x5D, 0x22, 0x34, 0x58, 0x76, 0x38, 0x36, 0x00, 0x5B, 0x24,
	0x07, 0x27, 0x56, 0x29, 0x7A, 0x02, 0x15, 0x2F, 0x44, 0x37, 0x1E, 0x1B,
	0x3E, 0x01, 0x09, 0x38, 0x0A, 0x26, 0x26, 0x2B, 0x25, 0x13, 0x3F, 0x26,
	0x18, 0x27, 0x55, 0x04, 0x31, 0x0E, 0x5E, 0x38, 0x3B, 0x11, 0x23, 0x2F,
	0x1B, 0x20, 0x18, 0x00, 0x47, 0x33, 0x09, 0x0C, 0x26, 0x1B, 0x29, 0x17,
	0x3D, 0x17, 0x2E, 0x4A, 0x2D, 0x18, 0x2A, 0x06, 0x17, 0x05, 0x29, 0x27,
	0x1A, 0x05, 0x2C, 0x22, 0x16, 0x43, 0x0C, 0x2D, 0x27, 0x6D, 0x22, 0x12,
	0x3F, 0x20, 0x1B, 0x38, 0x12, 0x02, 0x09, 0x21, 0x54, 0x18, 0x1A, 0x29,
	0x77, 0x02, 0x36, 0x2B, 0x58, 0x01, 0x19, 0x4A, 0x5A, 0x23, 0x17, 0x0B,
	0x51, 0x17, 0x28, 0x29, 0x27, 0x17, 0x1C, 0x1A, 0x71, 0x14, 0x2A, 0x17,
	0x3F, 0x36, 0x16, 0x31, 0x2A, 0x06, 0x2A, 0x5D, 0x2C, 0x17, 0x28, 0x24,
	0x26, 0x2E, 0x3D, 0x3A, 0x27, 0x21, 0x4A, 0x08, 0x44, 0x76, 0x27, 0x14,
	0x5B, 0x31, 0x75, 0x5E, 0x16, 0x58, 0x52, 0x03, 0x1D, 0x19, 0x21, 0x2A,
	0x2C, 0x2F, 0x27, 0x05, 0x18, 0x32, 0x05, 0x2B, 0x16, 0x03, 0x6D, 0x1B,
	0x3B, 0x38, 0x5E, 0x0F, 0x15, 0x2C, 0x2D, 0x2D, 0x7B, 0x1E, 0x0D, 0x1D,
	0x59, 0x0D, 0x5E, 0x0E, 0x07, 0x3B, 0x1B, 0x1F, 0x06, 0x38, 0x09, 0x1A,
	0x2D, 0x0D, 0x27, 0x29, 0x18, 0x2D, 0x02, 0x09, 0x0D, 0x35, 0x0A, 0x28,
	0x5F, 0x1C, 0x25, 0x59, 0x2A, 0x38, 0x31, 0x33, 0x06, 0x0E, 0x26, 0x26,
	0x28, 0x1B, 0x39, 0x17, 0x06, 0x0E, 0x47, 0x0F, 0x59, 0x13, 0x17, 0x23,
	0x23, 0x26, 0x59, 0x36, 0x35, 0x08, 0x5E, 0x18, 0x16, 0x2F, 0x4A, 0x26,
	0x1D, 0x27, 0x5F, 0x4A, 0x01, 0x25, 0x25, 0x1D, 0x50, 0x18, 0x1D, 0x06,
	0x15, 0x31, 0x5B, 0x0A, 0x33, 0x0A, 0x02, 0x5F, 0x00, 0x28, 0x43, 0x50,
	0x57, 0x19, 0x20, 0x2F, 0x30, 0x08, 0x1F, 0x20, 0x18, 0x37, 0x24, 0x3B,
	0x05, 0x1E, 0x29, 0x03, 0x0F, 0x15, 0x28, 0x50, 0x0B, 0x5D, 0x73, 0x35,
	0x2D, 0x41, 0x0A, 0x0A, 0x59, 0x36, 0x25, 0x11, 0x15, 0x3E, 0x06, 0x01,
	0x39, 0x29, 0x2B, 0x11, 0x28, 0x2F, 0x26, 0x0D, 0x3B, 0x27, 0x5F, 0x1A,
	0x3B, 0x56, 0x29, 0x5D, 0x18, 0x1F, 0x22, 0x26, 0x20, 0x24, 0x3D, 0x31,
	0x2B, 0x08, 0x04, 0x0B, 0x12, 0x38, 0x04, 0x32, 0x1E, 0x18, 0x14, 0x12,
	0x16, 0x0F, 0x33, 0x06, 0x0A, 0x70, 0x01, 0x19, 0x36, 0x1A, 0x74, 0x2B,
	0x2D, 0x34, 0x04, 0x33, 0x1B, 0x10, 0x2D, 0x00, 0x0F, 0x5D, 0x2E, 0x00,
	0x1F, 0x7A, 0x1E, 0x27, 0x1B, 0x2F, 0x2A, 0x00, 0x04, 0x07, 0x1D, 0x31,
	0x0D, 0x59, 0x0F, 0x1F, 0x74, 0x0E, 0x38, 0x02, 0x33, 0x16, 0x01, 0x28,
	0x06, 0x5E, 0x31, 0x04, 0x4E, 0x28, 0x59, 0x2C, 0x35, 0x17, 0x03, 0x04,
	0x09, 0x3B, 0x55, 0x29, 0x40, 0x08, 0x34, 0x2D, 0x38, 0x02, 0x3A, 0x36,
	0x24, 0x17, 0x13, 0x20, 0x1F, 0x03, 0x1E, 0x05, 0x6D, 0x1A, 0x2D, 0x02,
	0x1C, 0x23, 0x20, 0x27, 0x2D, 0x5D, 0x77, 0x09, 0x24, 0x02, 0x1C, 0x77,
	0x1A, 0x53, 0x08, 0x1B, 0x76, 0x00, 0x36, 0x1C, 0x3A, 0x0E, 0x36, 0x36,
	0x04, 0x2A, 0x24, 0x2F, 0x0D, 0x1C, 0x00, 0x77, 0x03, 0x12, 0x45, 0x53,
	0x12, 0x0E, 0x2F, 0x1F, 0x29, 0x2C, 0x05, 0x54, 0x23, 0x3D, 0x11, 0x1C,
	0x0D, 0x05, 0x1D, 0x04, 0x3A, 0x13, 0x03, 0x1C, 0x32, 0x00, 0x2A, 0x41,
	0x18, 0x2E, 0x05, 0x11, 0x22, 0x5A, 0x38, 0x3A, 0x12, 0x5B, 0x1B, 0x24,
	0x3F, 0x2D, 0x1A, 0x31, 0x2F, 0x21, 0x54, 0x00, 0x3A, 0x7B, 0x27, 0x31,
	0x3F, 0x44, 0x16, 0x09, 0x19, 0x2C, 0x40, 0x01, 0x25, 0x31, 0x37, 0x3A,
	0x27, 0x2E, 0x52, 0x5F, 0x32, 0x2E, 0x1B, 0x3B, 0x2A, 0x23, 0x1A, 0x5B,
	0x05, 0x04, 0x24, 0x2D, 0x22, 0x0A, 0x01, 0x09, 0x10, 0x14, 0x39, 0x07,
	0x32, 0x2E, 0x00, 0x55, 0x07, 0x5C, 0x30, 0x35, 0x34, 0x16, 0x31, 0x23,
	0x16, 0x24, 0x2C, 0x27, 0x2F, 0x0E, 0x2A, 0x02, 0x27, 0x0C, 0x02, 0x18,
	0x0D, 0x2D, 0x70, 0x08, 0x35, 0x1D, 0x04, 0x34, 0x20, 0x2E, 0x2C, 0x5D,
	0x36, 0x20, 0x52, 0x28, 0x01, 0x08, 0x1A, 0x12, 0x1C, 0x5C, 0x24, 0x26,
	0x4A, 0x07, 0x40, 0x04, 0x16, 0x03, 0x04, 0x38, 0x33, 0x2D, 0x02, 0x2A,
	0x1B, 0x2B, 0x08, 0x51, 0x45, 0x3B, 0x3B, 0x22, 0x00, 0x1E, 0x07, 0x29,
	0x01, 0x52, 0x28, 0x05, 0x37, 0x39, 0x10, 0x20, 0x24, 0x33, 0x2F, 0x10,
	0x3A, 0x13, 0x0B, 0x29, 0x36, 0x36, 0x52, 0x36, 0x2E, 0x0A, 0x2B, 0x1C,
	0x3A, 0x24, 0x07, 0x2B, 0x03, 0x70, 0x19, 0x37, 0x2C, 0x18, 0x0E, 0x3F,
	0x19, 0x1D, 0x29, 0x72, 0x3B, 0x14, 0x5B, 0x09, 0x2C, 0x34, 0x08, 0x5B,
	0x3A, 0x16, 0x3B, 0x2E, 0x17, 0x1A, 0x73, 0x2B, 0x1B, 0x3E, 0x5E, 0x0C,
	0x27, 0x04, 0x23, 0x1F, 0x11, 0x07, 0x27, 0x58, 0x52, 0x12, 0x23, 0x33,
	0x07, 0x52, 0x2D, 0x22, 0x28, 0x5F, 0x0F, 0x37, 0x22, 0x57, 0x1B, 0x3D,
	0x07, 0x02, 0x53, 0x08, 0x04, 0x0C, 0x01, 0x0A, 0x05, 0x3E, 0x10, 0x2F,
	0x24, 0x0C, 0x09, 0x2E, 0x0B, 0x57, 0x57, 0x3D, 0x09, 0x35, 0x09, 0x07,
	0x25, 0x27, 0x3F, 0x31, 0x5C, 0x38, 0x1B, 0x36, 0x57, 0x07, 0x39, 0x16,
	0x5D, 0x08, 0x58, 0x09, 0x12, 0x55, 0x4E, 0x56, 0x1F, 0x08, 0x2E, 0x4E,
	0x5E, 0x1E, 0x70, 0x5E, 0x03, 0x20, 0x07, 0x01, 0x3C, 0x36, 0x00, 0x13,
	0x72, 0x19, 0x22, 0x25, 0x3D, 0x24, 0x23, 0x17, 0x36, 0x29, 0x35, 0x1F,
	0x36, 0x22, 0x13, 0x29, 0x5E, 0x30, 0x1E, 0x5D, 0x09, 0x09, 0x36, 0x19,
	0x2D, 0x24, 0x36, 0x39, 0x27, 0x03, 0x32, 0x5E, 0x36, 0x09, 0x00, 0x07,
	0x0A, 0x39, 0x3B, 0x38, 0x74, 0x15, 0x4A, 0x38, 0x2A, 0x2D, 0x07, 0x03,
	0x5E, 0x29, 0x26, 0x5F, 0x15, 0x2F, 0x0F, 0x75, 0x3A, 0x4A, 0x28, 0x0C,
	0x3B, 0x22, 0x0D, 0x01, 0x01, 0x15, 0x0E, 0x30, 0x5F, 0x5D, 0x74, 0x34,
	0x27, 0x20, 0x38, 0x37, 0x3A, 0x0E, 0x21, 0x40, 0x11, 0x1C, 0x50, 0x29,
	0x40, 0x08, 0x0D, 0x30, 0x36, 0x06, 0x77, 0x1E, 0x38, 0x57, 0x29, 0x31,
	0x22, 0x34, 0x1C, 0x3F, 0x33, 0x5F, 0x26, 0x2A, 0x0D, 0x33, 0x0B, 0x2C,
	0x3A, 0x1B, 0x6D, 0x2E, 0x34, 0x1F, 0x3D, 0x33, 0x3B, 0x26, 0x14, 0x1B,
	0x34, 0x43, 0x03, 0x3D, 0x0E, 0x0D, 0x27, 0x08, 0x2C, 0x3C, 0x04, 0x0A,
	0x12, 0x38, 0x59, 0x0C, 0x0B, 0x51, 0x0F, 0x01, 0x10, 0x1E, 0x07, 0x05,
	0x02, 0x36, 0x21, 0x0E, 0x0C, 0x03, 0x18, 0x1C, 0x58, 0x23, 0x59, 0x21,
	0x23, 0x39, 0x3E, 0x24, 0x08, 0x36, 0x05, 0x0D, 0x59, 0x28, 0x5D, 0x1B,
	0x5F, 0x02, 0x1A, 0x08, 0x2C, 0x5C, 0x0F, 0x71, 0x34, 0x1B, 0x24, 0x11,
	0x77, 0x1D, 0x37, 0x0A, 0x1C, 0x23, 0x1D, 0x16, 0x1B, 0x0A, 0x3A, 0x23,
	0x17, 0x3D, 0x27, 0x2D, 0x24, 0x30, 0x5A, 0x1A, 0x77, 0x0F, 0x50, 0x1B,
	0x1E, 0x3A, 0x3A, 0x59, 0x27, 0x0C, 0x23, 0x55, 0x59, 0x0F, 0x0C, 0x6D,
	0x3B, 0x27, 0x0F, 0x05, 0x00, 0x47, 0x06, 0x1C, 0x07, 0x31, 0x26, 0x06,
	0x5C, 0x3C, 0x08, 0x09, 0x2C, 0x09, 0x13, 0x0B, 0x5B, 0x16, 0x19, 0x5B,
	0x3B, 0x1F, 0x27, 0x3F, 0x1A, 0x7A, 0x06, 0x0D, 0x0C, 0x3F, 0x08, 0x0D,
	0x0D, 0x39, 0x0C, 0x76, 0x3C, 0x54, 0x1E, 0x06, 0x77, 0x19, 0x4A, 0x3E,
	0x01, 0x29, 0x1A, 0x4E, 0x41, 0x0F, 0x04, 0x3F, 0x39, 0x3C, 0x07, 0x05,
	0x29, 0x07, 0x36, 0x32, 0x24, 0x25, 0x50, 0x5B, 0x5A, 0x16, 0x1F, 0x28,
	0x0B, 0x1E, 0x28, 0x43, 0x32, 0x08, 0x5A, 0x05, 0x23, 0x32, 0x41, 0x28,
	0x24, 0x1A, 0x56, 0x07, 0x39, 0x36, 0x47, 0x0B, 0x08, 0x3D, 0x38, 0x0E,
	0x2D, 0x2F, 0x44, 0x26, 0x05, 0x0A, 0x0F, 0x53, 0x27, 0x24, 0x2C, 0x14,
	0x27, 0x0F, 0x39, 0x51, 0x3B, 0x05, 0x12, 0x3D, 0x14, 0x1D, 0x58, 0x38,
	0x5C, 0x31, 0x3E, 0x21, 0x0B, 0x34, 0x32, 0x20, 0x1A, 0x77, 0x1C, 0x09,
	0x3E, 0x38, 0x38, 0x02, 0x4A, 0x1A, 0x32, 0x26, 0x1E, 0x11, 0x22, 0x05,
	0x18, 0x00, 0x03, 0x3A, 0x12, 0x0E, 0x1D, 0x10, 0x1C, 0x5F, 0x24, 0x01,
	0x16, 0x39, 0x33, 0x10, 0x06, 0x2F, 0x19, 0x58, 0x29, 0x5F, 0x26, 0x38,
	0x33, 0x12, 0x5D, 0x06, 0x0D, 0x5A, 0x2A, 0x1D, 0x19, 0x56, 0x3D, 0x27,
	0x55, 0x36, 0x3C, 0x33, 0x0C, 0x22, 0x13, 0x5F, 0x44, 0x09, 0x47, 0x0F,
	0x5E, 0x5D, 0x17, 0x09, 0x56, 0x39, 0x59, 0x10, 0x2D, 0x08, 0x5E, 0x5A,
	0x74, 0x03, 0x2C, 0x5E, 0x52, 0x0C, 0x1F, 0x51, 0x16, 0x3A, 0x77, 0x39,
	0x4A, 0x1B, 0x21, 0x25, 0x38, 0x09, 0x08, 0x19, 0x2F, 0x2B, 0x2A, 0x5B,
	0x23, 0x0E, 0x3D, 0x00, 0x04, 0x31, 0x25, 0x02, 0x11, 0x3A, 0x1B, 0x0C,
	0x24, 0x16, 0x3A, 0x39, 0x24, 0x2A, 0x2B, 0x1A, 0x07, 0x7B, 0x39, 0x0A,
	0x29, 0x3D, 0x26, 0x27, 0x55, 0x1F, 0x40, 0x32, 0x06, 0x0E, 0x1E, 0x32,
	0x11, 0x1B, 0x04, 0x57, 0x0A, 0x32, 0x0D, 0x0D, 0x20, 0x0C, 0x36, 0x0E,
	0x28, 0x39, 0x05, 0x33, 0x59, 0x38, 0x5F, 0x40, 0x6D, 0x1C, 0x57, 0x05,
	0x3E, 0x05, 0x3C, 0x10, 0x38, 0x53, 0x05, 0x3F, 0x2C, 0x28, 0x5C, 0x06,
	0x01, 0x32, 0x02, 0x19, 0x2B, 0x02, 0x27, 0x1E, 0x0C, 0x09, 0x3B, 0x00,
	0x3E, 0x29, 0x0D, 0x1C, 0x30, 0x02, 0x58, 0x72, 0x05, 0x51, 0x1E, 0x0A,
	0x2F, 0x39, 0x54, 0x1F, 0x27, 0x0C, 0x0E, 0x57, 0x22, 0x52, 0x04, 0x5E,
	0x58, 0x3B, 0x2A, 0x26, 0x06, 0x18, 0x24, 0x1E, 0x24, 0x5E, 0x2E, 0x02,
	0x12, 0x15, 0x0F, 0x51, 0x2B, 0x0C, 0x27, 0x24, 0x19, 0x0D, 0x39, 0x35,
	0x0A, 0x54, 0x3C, 0x1D, 0x0C, 0x34, 0x2E, 0x5E, 0x3B, 0x7A, 0x1C, 0x13,
	0x03, 0x3B, 0x26, 0x2B, 0x30, 0x29, 0x40, 0x14, 0x36, 0x0F, 0x2D, 0x12,
	0x7B, 0x05, 0x2D, 0x5C, 0x1E, 0x69, 0x00, 0x29, 0x3A, 0x5D, 0x2D, 0x3F,
	0x2E, 0x3C, 0x21, 0x2A, 0x3B, 0x35, 0x5F, 0x59, 0x32, 0x38, 0x54, 0x59,
	0x3D, 0x36, 0x2D, 0x07, 0x16, 0x05, 0x16, 0x55, 0x0C, 0x07, 0x1B, 0x21,
	0x3A, 0x0C, 0x1C, 0x13, 0x69, 0x1B, 0x0F, 0x3B, 0x25, 0x0D, 0x0D, 0x53,
	0x34, 0x5E, 0x29, 0x27, 0x2A, 0x5D, 0x27, 0x34, 0x03, 0x17, 0x1F, 0x1C,
	0x16, 0x26, 0x11, 0x16, 0x0E, 0x04, 0x1D, 0x0E, 0x5E, 0x01, 0x34, 0x26,
	0x17, 0x1C, 0x3C, 0x69, 0x1D, 0x0E, 0x0A, 0x23, 0x03, 0x58, 0x50, 0x5C,
	0x07, 0x21, 0x08, 0x57, 0x1A, 0x3E, 0x32, 0x0A, 0x19, 0x41, 0x5A, 0x28,
	0x18, 0x34, 0x04, 0x58, 0x30, 0x58, 0x56, 0x2F, 0x05, 0x06, 0x5B, 0x29,
	0x05, 0x3D, 0x10, 0x3B, 0x24, 0x1A, 0x5A, 0x01, 0x05, 0x33, 0x04, 0x2F,
	0x0D, 0x1D, 0x58, 0x06, 0x06, 0x75, 0x36, 0x0A, 0x02, 0x40, 0x2A, 0x2D,
	0x38, 0x1E, 0x5A, 0x20, 0x55, 0x30, 0x59, 0x23, 0x18, 0x2F, 0x0D, 0x59,
	0x1D, 0x7B, 0x22, 0x15, 0x5E, 0x08, 0x6D, 0x5A, 0x18, 0x04, 0x3F, 0x00,
	0x3B, 0x54, 0x2D, 0x0D, 0x31, 0x38, 0x1B, 0x57, 0x2E, 0x28, 0x34, 0x07,
	0x58, 0x3C, 0x37, 0x14, 0x55, 0x2B, 0x29, 0x1B, 0x0E, 0x2F, 0x1E, 0x1E,
	0x2D, 0x3A, 0x54, 0x04, 0x09, 0x3B, 0x23, 0x2E, 0x29, 0x11, 0x14, 0x0E,
	0x23, 0x04, 0x39, 0x13, 0x14, 0x54, 0x27, 0x2D, 0x77, 0x0F, 0x11, 0x09,
	0x21, 0x15, 0x1D, 0x51, 0x20, 0x2D, 0x0C, 0x0F, 0x57, 0x3C, 0x18, 0x0D,
	0x2B, 0x0D, 0x17, 0x0F, 0x21, 0x0E, 0x22, 0x16, 0x26, 0x17, 0x14, 0x0C,
	0x5F, 0x5A, 0x20, 0x07, 0x31, 0x08, 0x3F, 0x77, 0x3F, 0x34, 0x58, 0x05,
	0x2F, 0x5D, 0x27, 0x08, 0x21, 0x69, 0x20, 0x17, 0x5A, 0x00, 0x38, 0x2E,
	0x53, 0x06, 0x5D, 0x2B, 0x34, 0x13, 0x57, 0x39, 0x24, 0x5B, 0x50, 0x58,
	0x2E, 0x0C, 0x3B, 0x2A, 0x5E, 0x32, 0x06, 0x47, 0x33, 0x37, 0x53, 0x05,
	0x08, 0x02, 0x3E, 0x1B, 0x74, 0x2A, 0x29, 0x2C, 0x05, 0x20, 0x5B, 0x0A,
	0x24, 0x11, 0x73, 0x29, 0x10, 0x26, 0x3B, 0x16, 0x36, 0x4E, 0x34, 0x1E,
	0x28, 0x39, 0x19, 0x01, 0x39, 0x7B, 0x1C, 0x53, 0x08, 0x52, 0x70, 0x27,
	0x52, 0x5E, 0x01, 0x13, 0x5A, 0x2F, 0x5C, 0x0C, 0x06, 0x2D, 0x39, 0x5D,
	0x11, 0x72, 0x3C, 0x27, 0x38, 0x01, 0x71, 0x20, 0x04, 0x1F, 0x0C, 0x70,
	0x47, 0x06, 0x38, 0x5A, 0x2D, 0x55, 0x38, 0x09, 0x12, 0x3B, 0x02, 0x15,
	0x08, 0x24, 0x2D, 0x28, 0x57, 0x3B, 0x3A, 0x07, 0x0A, 0x02, 0x20, 0x40,
	0x34, 0x47, 0x30, 0x36, 0x3B, 0x26, 0x2E, 0x03, 0x5D, 0x0A, 0x2A, 0x5B,
	0x36, 0x25, 0x07, 0x23, 0x1E, 0x2F, 0x3A, 0x38, 0x76, 0x39, 0x51, 0x18,
	0x19, 0x21, 0x1B, 0x17, 0x09, 0x3C, 0x74, 0x06, 0x36, 0x06, 0x11, 0x15,
	0x19, 0x33, 0x3A, 0x1A, 0x20, 0x0D, 0x33, 0x18, 0x21, 0x34, 0x5E, 0x2B,
	0x3C, 0x5A, 0x2B, 0x06, 0x29, 0x3B, 0x18, 0x20, 0x3F, 0x31, 0x0D, 0x07,
	0x6D, 0x1C, 0x2C, 0x38, 0x22, 0x27, 0x5A, 0x00, 0x08, 0x18, 0x29, 0x5C,
	0x55, 0x29, 0x25, 0x0D, 0x39, 0x58, 0x37, 0x58, 0x23, 0x0E, 0x0E, 0x18,
	0x1D, 0x35, 0x2B, 0x15, 0x04, 0x31, 0x33, 0x54, 0x23, 0x39, 0x28, 0x25,
	0x01, 0x03, 0x59, 0x02, 0x15, 0x02, 0x26, 0x14, 0x5D, 0x06, 0x20, 0x53,
	0x0A, 0x1A, 0x2E, 0x5F, 0x10, 0x37, 0x0F, 0x34, 0x3E, 0x16, 0x3E, 0x1A,
	0x0B, 0x55, 0x11, 0x3E, 0x5A, 0x33, 0x27, 0x39, 0x5D, 0x12, 0x20, 0x5B,
	0x34, 0x0B, 0x00, 0x24, 0x5C, 0x50, 0x20, 0x09, 0x36, 0x3B, 0x2A, 0x39,
	0x3F, 0x21, 0x36, 0x4E, 0x0C, 0x25, 0x26, 0x26, 0x0C, 0x34, 0x3E, 0x05,
	0x3B, 0x2E, 0x02, 0x06, 0x11, 0x0D, 0x06, 0x45, 0x19, 0x0A, 0x55, 0x39,
	0x0C, 0x5A, 0x08, 0x1A, 0x29, 0x3B, 0x11, 0x0A, 0x3F, 0x2F, 0x29, 0x04,
	0x03, 0x06, 0x2E, 0x09, 0x31, 0x7A, 0x59, 0x28, 0x02, 0x2D, 0x70, 0x0B,
	0x31, 0x58, 0x2C, 0x73, 0x5D, 0x20, 0x02, 0x1E, 0x7A, 0x2F, 0x06, 0x22,
	0x40, 0x35, 0x0F, 0x35, 0x04, 0x29, 0x2B, 0x39, 0x57, 0x1A, 0x11, 0x13,
	0x1E, 0x0C, 0x41, 0x26, 0x14, 0x06, 0x31, 0x58, 0x5A, 0x2D, 0x5F, 0x04,
	0x57, 0x2F, 0x2D, 0x2E, 0x17, 0x3C, 0x3A, 0x3B, 0x38, 0x12, 0x03, 0x11,
	0x2D, 0x2B, 0x54, 0x22, 0x04, 0x3B, 0x5A, 0x2A, 0x57, 0x25, 0x37, 0x05,
	0x2E, 0x5C, 0x3D, 0x2E, 0x07, 0x07, 0x19, 0x38, 0x0C, 0x0A, 0x33, 0x36,
	0x04, 0x0B, 0x09, 0x13, 0x5E, 0x20, 0x37, 0x3F, 0x06, 0x57, 0x1A, 0x7A,
	0x38, 0x25, 0x27, 0x20, 0x7B, 0x26, 0x25, 0x1A, 0x2F, 0x17, 0x02, 0x33,
	0x06, 0x11, 0x3B, 0x3B, 0x35, 0x3C, 0x00, 0x36, 0x22, 0x0E, 0x1C, 0x09,
	0x73, 0x3B, 0x2A, 0x1C, 0x24, 0x2F, 0x15, 0x07, 0x01, 0x2D, 0x35, 0x22,
	0x57, 0x20, 0x2D, 0x20, 0x2A, 0x07, 0x5F, 0x1E, 0x05, 0x0D, 0x0A, 0x25,
	0x13, 0x03, 0x1B, 0x24, 0x08, 0x04, 0x11, 0x2E, 0x12, 0x20, 0x22, 0x6D,
	0x29, 0x23, 0x18, 0x3D, 0x70, 0x21, 0x05, 0x5C, 0x18, 0x20, 0x59, 0x16,
	0x21, 0x12, 0x08, 0x2F, 0x50, 0x0B, 0x05, 0x77, 0x03, 0x16, 0x0C, 0x2D,
	0x12, 0x01, 0x37, 0x0A, 0x1F, 0x6D, 0x39, 0x29, 0x1C, 0x32, 0x24, 0x5C,
	0x33, 0x5E, 0x08, 0x1B, 0x5B, 0x0B, 0x1D, 0x31, 0x34, 0x19, 0x13, 0x16,
	0x1E, 0x0E, 0x19, 0x0E, 0x3E, 0x1B, 0x01, 0x00, 0x0A, 0x0A, 0x3E, 0x24,
	0x5A, 0x2C, 0x1B, 0x00, 0x71, 0x5C, 0x55, 0x06, 0x1B, 0x1A, 0x0D, 0x13,
	0x28, 0x0F, 0x23, 0x16, 0x0D, 0x0C, 0x01, 0x10, 0x18, 0x4A, 0x0C, 0x3F,
	0x0F, 0x2A, 0x52, 0x03, 0x12, 0x76, 0x43, 0x00, 0x2B, 0x39, 0x29, 0x14,
	0x54, 0x3B, 0x21, 0x24, 0x1C, 0x34, 0x39, 0x0D, 0x09, 0x3E, 0x54, 0x3F,
	0x39, 0x15, 0x5E, 0x32, 0x00, 0x01, 0x6D, 0x39, 0x00, 0x2C, 0x00, 0x0C,
	0x3D, 0x57, 0x21, 0x02, 0x3B, 0x3E, 0x38, 0x0C, 0x58, 0x23, 0x03, 0x00,
	0x2D, 0x0C, 0x0F, 0x18, 0x54, 0x08, 0x1F, 0x17, 0x3A, 0x25, 0x56, 0x19,
	0x32, 0x59, 0x53, 0x02, 0x2D, 0x08, 0x00, 0x19, 0x36, 0x12, 0x2C, 0x3E,
	0x2C, 0x28, 0x2C, 0x09, 0x00, 0x20, 0x0A, 0x44, 0x15, 0x26, 0x54, 0x45,
	0x3C, 0x17, 0x2A, 0x11, 0x09, 0x39, 0x09, 0x36, 0x20, 0x41, 0x23, 0x72,
	0x5B, 0x0E, 0x25, 0x5D, 0x26, 0x24, 0x2B, 0x0A, 0x3B, 0x21, 0x0E, 0x37,
	0x3F, 0x26, 0x34, 0x5A, 0x06, 0x58, 0x25, 0x07, 0x29, 0x16, 0x38, 0x26,
	0x0A, 0x3F, 0x14, 0x21, 0x1A, 0x20, 0x23, 0x13, 0x2F, 0x0E, 0x1B, 0x47,
	0x27, 0x39, 0x00, 0x23, 0x28, 0x0D, 0x3F, 0x3E, 0x69, 0x0F, 0x37, 0x26,
	0x5B, 0x3B, 0x55, 0x37, 0x59, 0x5A, 0x75, 0x59, 0x2C, 0x1F, 0x5A, 0x35,
	0x07, 0x56, 0x1C, 0x58, 0x73, 0x06, 0x25, 0x5D, 0x3F, 0x2C, 0x19, 0x09,
	0x34, 0x22, 0x00, 0x0D, 0x06, 0x22, 0x38, 0x37, 0x24, 0x13, 0x5A, 0x1C,
	0x70, 0x0A, 0x30, 0x5F, 0x00, 0x25, 0x5A, 0x08, 0x08, 0x1F, 0x26, 0x55,
	0x1B, 0x37, 0x5D, 0x70, 0x1F, 0x09, 0x5D, 0x07, 0x30, 0x38, 0x25, 0x1A,
	0x39, 0x0F, 0x07, 0x39, 0x34, 0x08, 0x36, 0x28, 0x15, 0x58, 0x27, 0x10,
	0x3D, 0x36, 0x3E, 0x09, 0x1A, 0x29, 0x2D, 0x28, 0x3E, 0x73, 0x14, 0x27,
	0x17, 0x0C, 0x72, 0x0D, 0x29, 0x25, 0x05, 0x13, 0x26, 0x0E, 0x19, 0x44,
	0x0C, 0x08, 0x07, 0x20, 0x25, 0x35, 0x1C, 0x2A, 0x0C, 0x27, 0x37, 0x35,
	0x52, 0x1B, 0x52, 0x2D, 0x3F, 0x2A, 0x1A, 0x0F, 0x3B, 0x2B, 0x55, 0x1F,
	0x1B, 0x70, 0x36, 0x32, 0x57, 0x19, 0x24, 0x34, 0x31, 0x34, 0x12, 0x75,
	0x00, 0x34, 0x1F, 0x44, 0x75, 0x2F, 0x25, 0x28, 0x05, 0x7B, 0x07, 0x00,
	0x3E, 0x2C, 0x76, 0x1A, 0x34, 0x0C, 0x5A, 0x24, 0x02, 0x34, 0x24, 0x25,
	0x10, 0x02, 0x22, 0x1C, 0x1C, 0x31, 0x1C, 0x27, 0x58, 0x39, 0x28, 0x58,
	0x29, 0x1B, 0x1A, 0x36, 0x1D, 0x25, 0x57, 0x1F, 0x08, 0x25, 0x37, 0x1D,
	0x05, 0x04, 0x47, 0x15, 0x24, 0x2F, 0x2F, 0x0B, 0x16, 0x26, 0x25, 0x14,
	0x1B, 0x03, 0x04, 0x20, 0x13, 0x0E, 0x22, 0x09, 0x33, 0x23, 0x01, 0x36,
	0x3F, 0x5C, 0x72, 0x14, 0x2A, 0x04, 0x23, 0x6D, 0x09, 0x29, 0x23, 0x3A,
	0x1A, 0x39, 0x58, 0x07, 0x08, 0x75, 0x03, 0x38, 0x25, 0x5F, 0x27, 0x00,
	0x22, 0x03, 0x1E, 0x15, 0x20, 0x2A, 0x18, 0x39, 0x2B, 0x21, 0x09, 0x03,
	0x19, 0x0B, 0x06, 0x55, 0x1A, 0x08, 0x27, 0x2D, 0x15, 0x3C, 0x06, 0x21,
	0x38, 0x13, 0x34, 0x0A, 0x12, 0x20, 0x50, 0x0A, 0x19, 0x73, 0x35, 0x53,
	0x06, 0x1A, 0x13, 0x1E, 0x11, 0x03, 0x52, 0x2F, 0x2A, 0x58, 0x14, 0x5E,
	0x34, 0x3F, 0x0D, 0x41, 0x5A, 0x3A, 0x19, 0x58, 0x06, 0x04, 0x20, 0x5D,
	0x07, 0x57, 0x08, 0x0F, 0x1E, 0x57, 0x22, 0x44, 0x30, 0x00, 0x10, 0x16,
	0x21, 0x05, 0x05, 0x35, 0x00, 0x0F, 0x30, 0x14, 0x03, 0x57, 0x59, 0x26,
	0x43, 0x1B, 0x3C, 0x11, 0x16, 0x19, 0x04, 0x41, 0x11, 0x18, 0x5B, 0x37,
	0x56, 0x3C, 0x7B, 0x5A, 0x14, 0x02, 0x09, 0x24, 0x1A, 0x11, 0x21, 0x22,
	0x2F, 0x1A, 0x51, 0x5E, 0x3C, 0x03, 0x59, 0x37, 0x59, 0x2E, 0x37, 0x43,
	0x59, 0x17, 0x2A, 0x0B, 0x22, 0x58, 0x00, 0x3B, 0x33, 0x15, 0x0E, 0x22,
	0x53, 0x21, 0x38, 0x25, 0x3E, 0x31, 0x04, 0x1F, 0x24, 0x2A, 0x32, 0x31,
	0x2F, 0x0E, 0x21, 0x18, 0x74, 0x55, 0x34, 0x1D, 0x04, 0x11, 0x25, 0x56,
	0x0D, 0x01, 0x1B, 0x0B, 0x53, 0x34, 0x0C, 0x14, 0x20, 0x37, 0x18, 0x59,
	0x12, 0x29, 0x59, 0x38, 0x40, 0x2F, 0x02, 0x55, 0x38, 0x3B, 0x32, 0x59,
	0x33, 0x25, 0x38, 0x1B, 0x25, 0x04, 0x27, 0x5C, 0x31, 0x29, 0x18, 0x0A,
	0x5C, 0x28, 0x25, 0x08, 0x1E, 0x3D, 0x29, 0x25, 0x57, 0x57, 0x39, 0x17,
	0x5F, 0x33, 0x1C, 0x23, 0x24, 0x47, 0x06, 0x04, 0x53, 0x2E, 0x08, 0x0C,
	0x5F, 0x5B, 0x07, 0x36, 0x0B, 0x59, 0x58, 0x36, 0x1A, 0x0B, 0x59, 0x1A,
	0x1B, 0x23, 0x3B, 0x2D, 0x58, 0x0C, 0x2B, 0x11, 0x3D, 0x59, 0x0B, 0x38,
	0x3B, 0x37, 0x26, 0x15, 0x23, 0x27, 0x5B, 0x31, 0x14, 0x0F, 0x50, 0x1C,
	0x3F, 0x10, 0x59, 0x51, 0x0C, 0x27, 0x75, 0x0D, 0x04, 0x36, 0x1A, 0x74,
	0x0D, 0x0A, 0x01, 0x20, 0x31, 0x1F, 0x0C, 0x0A, 0x03, 0x2C, 0x3D, 0x2C,
	0x36, 0x59, 0x26, 0x16, 0x52, 0x2D, 0x1B, 0x0D, 0x02, 0x53, 0x02, 0x44,
	0x77, 0x35, 0x14, 0x1E, 0x3B, 0x75, 0x25, 0x19, 0x1F, 0x29, 0x35, 0x0D,
	0x58, 0x34, 0x22, 0x28, 0x1F, 0x06, 0x3B, 0x01, 0x31, 0x04, 0x52, 0x1F,
	0x44, 0x24, 0x29, 0x20, 0x36, 0x33, 0x3A, 0x20, 0x11, 0x36, 0x52, 0x0E,
	0x1F, 0x39, 0x57, 0x5D, 0x14, 0x58, 0x13, 0x1E, 0x12, 0x7A, 0x14, 0x2E,
	0x2F, 0x33, 0x15, 0x04, 0x36, 0x39, 0x06, 0x1A, 0x03, 0x1B, 0x1D, 0x02,
	0x2A, 0x1A, 0x55, 0x25, 0x2C, 0x13, 0x43, 0x23, 0x01, 0x29, 0x29, 0x09,
	0x07, 0x1E, 0x12, 0x0B, 0x26, 0x58, 0x24, 0x3C, 0x33, 0x16, 0x06, 0x23,
	0x2A, 0x11, 0x3F, 0x04, 0x1C, 0x18, 0x28, 0x25, 0x55, 0x1A, 0x2E, 0x29,
	0x55, 0x24, 0x20, 0x2C, 0x27, 0x14, 0x13, 0x0C, 0x2D, 0x24, 0x35, 0x30,
	0x25, 0x1A, 0x16, 0x39, 0x0C, 0x09, 0x58, 0x73, 0x35, 0x58, 0x0C, 0x07,
	0x00, 0x03, 0x0E, 0x5E, 0x3D, 0x10, 0x0B, 0x0D, 0x5E, 0x3B, 0x2F, 0x2F,
	0x4E, 0x22, 0x23, 0x2D, 0x2D, 0x54, 0x2D, 0x52, 0x12, 0x34, 0x2C, 0x2B,
	0x20, 0x23, 0x3A, 0x37, 0x45, 0x2D, 0x0D, 0x35, 0x57, 0x5D, 0x3C, 0x77,
	0x1F, 0x14, 0x5C, 0x5D, 0x75, 0x06, 0x0F, 0x02, 0x01, 0x04, 0x05, 0x09,
	0x3B, 0x39, 0x0E, 0x5D, 0x33, 0x02, 0x3A, 0x33, 0x5D, 0x06, 0x1B, 0x2F,
	0x08, 0x0A, 0x26, 0x1C, 0x0E, 0x2A, 0x22, 0x00, 0x21, 0x59, 0x30, 0x29,
	0x17, 0x0F, 0x19, 0x37, 0x3E, 0x05, 0x16, 0x58, 0x03, 0x01, 0x53, 0x05,
	0x1A, 0x10, 0x55, 0x37, 0x2B, 0x44, 0x05, 0x3E, 0x35, 0x39, 0x0D, 0x10,
	0x16, 0x11, 0x3C, 0x01, 0x70, 0x1B, 0x0C, 0x0D, 0x1B, 0x35, 0x07, 0x2F,
	0x21, 0x5E, 0x3B, 0x5D, 0x38, 0x00, 0x58, 0x1B, 0x08, 0x0B, 0x00, 0x59,
	0x21, 0x26, 0x34, 0x2D, 0x5E, 0x0F, 0x22, 0x39, 0x5E, 0x18, 0x77, 0x22,
	0x03, 0x5C, 0x0A, 0x2D, 0x39, 0x06, 0x5B, 0x05, 0x33, 0x0E, 0x4A, 0x26,
	0x02, 0x13, 0x09, 0x02, 0x2B, 0x08, 0x36, 0x01, 0x2D, 0x01, 0x5E, 0x05,
	0x2E, 0x53, 0x17, 0x1D, 0x21, 0x5B, 0x37, 0x5E, 0x26, 0x2C, 0x00, 0x03,
	0x59, 0x08, 0x2D, 0x2B, 0x02, 0x1C, 0x2C, 0x2D, 0x15, 0x00, 0x20, 0x1B,
	0x0F, 0x27, 0x04, 0x22, 0x2C, 0x70, 0x3E, 0x28, 0x3B, 0x27, 0x21, 0x20,
	0x14, 0x01, 0x3B, 0x0D, 0x3A, 0x51, 0x1D, 0x5D, 0x2D, 0x03, 0x10, 0x19,
	0x06, 0x32, 0x58, 0x55, 0x07, 0x06, 0x2A, 0x21, 0x50, 0x5C, 0x1C, 0x70,
	0x04, 0x12, 0x19, 0x5F, 0x0B, 0x2B, 0x51, 0x5E, 0x02, 0x28, 0x16, 0x2B,
	0x36, 0x00, 0x08, 0x23, 0x24, 0x2B, 0x58, 0x16, 0x59, 0x18, 0x1A, 0x26,
	0x38, 0x1F, 0x57, 0x04, 0x0A, 0x74, 0x2F, 0x27, 0x3D, 0x0F, 0x21, 0x47,
	0x14, 0x1F, 0x1F, 0x16, 0x2D, 0x18, 0x21, 0x03, 0x2C, 0x1C, 0x1B, 0x1D,
	0x29, 0x18, 0x1E, 0x39, 0x34, 0x28, 0x69, 0x03, 0x27, 0x58, 0x06, 0x20,
	0x04, 0x35, 0x17, 0x27, 0x15, 0x1C, 0x16, 0x41, 0x0A, 0x77, 0x22, 0x07,
	0x0D, 0x3E, 0x10, 0x0D, 0x0B, 0x34, 0x13, 0x24, 0x01, 0x12, 0x58, 0x0F,
	0x34, 0x14, 0x33, 0x0C, 0x44, 0x21, 0x07, 0x37, 0x0A, 0x23, 0x21, 0x0F,
	0x22, 0x2A, 0x08, 0x0A, 0x1A, 0x2C, 0x0D, 0x58, 0x09, 0x18, 0x08, 0x5B,
	0x1D, 0x14, 0x34, 0x17, 0x3A, 0x5C, 0x7A, 0x3A, 0x2A, 0x3C, 0x38, 0x74,
	0x29, 0x12, 0x5D, 0x02, 0x7A, 0x0F, 0x3B, 0x19, 0x3C, 0x0F, 0x27, 0x58,
	0x37, 0x3F, 0x69, 0x1E, 0x13, 0x0F, 0x22, 0x2C, 0x38, 0x36, 0x0F, 0x0A,
	0x03, 0x19, 0x2E, 0x29, 0x05, 0x23, 0x07, 0x2D, 0x1F, 0x40, 0x12, 0x3B,
	0x12, 0x00, 0x19, 0x21, 0x34, 0x24, 0x3A, 0x3B, 0x30, 0x1F, 0x19, 0x56,
	0x5A, 0x2C, 0x2F, 0x53, 0x45, 0x05, 0x69, 0x0B, 0x3B, 0x07, 0x1B, 0x2C,
	0x00, 0x2E, 0x07, 0x19, 0x7A, 0x3C, 0x4A, 0x0C, 0x2A, 0x20, 0x23, 0x32,
	0x20, 0x38, 0x76, 0x0A, 0x53, 0x25, 0x3E, 0x6D, 0x0D, 0x02, 0x28, 0x2E,
	0x07, 0x2E, 0x16, 0x2B, 0x25, 0x1B, 0x3A, 0x18, 0x3C, 0x1B, 0x38, 0x19,
	0x31, 0x0C, 0x27, 0x69, 0x1D, 0x34, 0x3D, 0x1E, 0x2E, 0x38, 0x08, 0x2D,
	0x09, 0x0C, 0x5B, 0x30, 0x23, 0x2E, 0x1B, 0x1E, 0x19, 0x27, 0x2F, 0x12,
	0x39, 0x2B, 0x16, 0x00, 0x15, 0x14, 0x0E, 0x41, 0x1A, 0x30, 0x0F, 0x57,
	0x17, 0x18, 0x71, 0x34, 0x4A, 0x0F, 0x5D, 0x33, 0x25, 0x37, 0x03, 0x5A,
	0x77, 0x55, 0x0C, 0x07, 0x04, 0x21, 0x21, 0x31, 0x17, 0x00, 0x7A, 0x55,
	0x56, 0x5C, 0x1F, 0x2C, 0x22, 0x00, 0x2C, 0x5E, 0x36, 0x55, 0x51, 0x5E,
	0x01, 0x36, 0x29, 0x0E, 0x2A, 0x5D, 0x13, 0x2F, 0x28, 0x28, 0x00, 0x24,
	0x1D, 0x10, 0x36, 0x3F, 0x09, 0x03, 0x13, 0x29, 0x3B, 0x70, 0x3A, 0x0D,
	0x17, 0x1B, 0x77, 0x15, 0x34, 0x27, 0x53, 0x0A, 0x3E, 0x13, 0x05, 0x00,
	0x2B, 0x43, 0x27, 0x05, 0x11, 0x11, 0x55, 0x51, 0x5B, 0x26, 0x26, 0x1B,
	0x20, 0x5E, 0x05, 0x0C, 0x35, 0x0E, 0x05, 0x3E, 0x76, 0x0F, 0x0B, 0x17,
	0x20, 0x2B, 0x5A, 0x08, 0x1C, 0x24, 0x18, 0x3E, 0x54, 0x20, 0x03, 0x13,
	0x36, 0x2F, 0x57, 0x08, 0x69, 0x09, 0x06, 0x5E, 0x1F, 0x29, 0x20, 0x58,
	0x2F, 0x2F, 0x33, 0x3D, 0x16, 0x25, 0x33, 0x31, 0x09, 0x35, 0x27, 0x05,
	0x17, 0x1B, 0x26, 0x0C, 0x0C, 0x30, 0x3F, 0x00, 0x57, 0x2A, 0x23, 0x20,
	0x0E, 0x5D, 0x53, 0x13, 0x5A, 0x16, 0x1B, 0x3B, 0x0E, 0x29, 0x06, 0x14,
	0x3A, 0x18, 0x19, 0x57, 0x19, 0x06, 0x01, 0x59, 0x05, 0x17, 0x3A, 0x77,
	0x22, 0x55, 0x0F, 0x04, 0x2D, 0x0B, 0x0C, 0x04, 0x3B, 0x05, 0x47, 0x19,
	0x3B, 0x01, 0x15, 0x09, 0x0A, 0x0B, 0x11, 0x21, 0x3D, 0x19, 0x38, 0x38,
	0x0D, 0x28, 0x16, 0x3A, 0x08, 0x28, 0x15, 0x2B, 0x24, 0x1E, 0x2E, 0x25,
	0x35, 0x3B, 0x0E, 0x28, 0x55, 0x0F, 0x24, 0x5D, 0x26, 0x0A, 0x33, 0x24,
	0x06, 0x36, 0x3A, 0x08, 0x21, 0x5D, 0x33, 0x1B, 0x12, 0x02, 0x32, 0x69,
	0x27, 0x17, 0x1D, 0x0F, 0x15, 0x3E, 0x50, 0x27, 0x29, 0x17, 0x24, 0x31,
	0x39, 0x5E, 0x38, 0x16, 0x59, 0x23, 0x0C, 0x0B, 0x1D, 0x0C, 0x57, 0x26,
	0x28, 0x3E, 0x0F, 0x04, 0x0A, 0x31, 0x0E, 0x59, 0x2B, 0x2D, 0x34, 0x2F,
	0x27, 0x1F, 0x06, 0x2C, 0x3F, 0x0A, 0x3A, 0x06, 0x38, 0x58, 0x1B, 0x05,
	0x22, 0x00, 0x26, 0x11, 0x0F, 0x0D, 0x2F, 0x01, 0x17, 0x00, 0x32, 0x21,
	0x22, 0x35, 0x16, 0x28, 0x3B, 0x59, 0x0C, 0x07, 0x2C, 0x76, 0x43, 0x18,
	0x2F, 0x18, 0x33, 0x22, 0x04, 0x03, 0x11, 0x7A, 0x0E, 0x15, 0x5E, 0x3D,
	0x14, 0x20, 0x02, 0x3F, 0x01, 0x11, 0x2F, 0x28, 0x21, 0x0F, 0x0B, 0x3A,
	0x19, 0x08, 0x0D, 0x17, 0x3A, 0x53, 0x3C, 0x0F, 0x75, 0x28, 0x17, 0x3A,
	0x23, 0x23, 0x58, 0x52, 0x23, 0x5F, 0x2E, 0x2F, 0x12, 0x29, 0x5F, 0x26,
	0x5B, 0x04, 0x21, 0x1B, 0x26, 0x3A, 0x00, 0x0B, 0x03, 0x17, 0x0E, 0x14,
	0x23, 0x40, 0x38, 0x35, 0x2A, 0x39, 0x18, 0x17, 0x35, 0x0E, 0x0B, 0x25,
	0x77, 0x04, 0x1B, 0x41, 0x38, 0x15, 0x5E, 0x16, 0x25, 0x3C, 0x0B, 0x06,
	0x08, 0x5E, 0x24, 0x27, 0x24, 0x2D, 0x09, 0x0A, 0x73, 0x02, 0x56, 0x2A,
	0x20, 0x0E, 0x08, 0x0B, 0x00, 0x2D, 0x3B, 0x23, 0x55, 0x18, 0x1F, 0x0F,
	0x36, 0x2E, 0x34, 0x06, 0x1A, 0x25, 0x2A, 0x00, 0x3A, 0x77, 0x5F, 0x16,
	0x5B, 0x18, 0x0E, 0x5E, 0x18, 0x41, 0x21, 0x24, 0x2E, 0x50, 0x39, 0x25,
	0x72, 0x27, 0x18, 0x41, 0x31, 0x31, 0x43, 0x0B, 0x0A, 0x09, 0x15, 0x39,
	0x23, 0x19, 0x5F, 0x20, 0x2B, 0x58, 0x28, 0x39, 0x75, 0x54, 0x09, 0x20,
	0x3E, 0x76, 0x1A, 0x03, 0x03, 0x0E, 0x2F, 0x22, 0x1B, 0x0F, 0x31, 0x21,
	0x04, 0x2C, 0x2A, 0x1B, 0x21, 0x19, 0x2D, 0x1F, 0x0D, 0x26, 0x34, 0x1B,
	0x18, 0x33, 0x0E, 0x25, 0x18, 0x19, 0x58, 0x72, 0x09, 0x15, 0x24, 0x27,
	0x0E, 0x2D, 0x11, 0x22, 0x5E, 0x0B, 0x22, 0x16, 0x25, 0x25, 0x3A, 0x3D,
	0x1B, 0x0B, 0x00, 0x74, 0x16, 0x55, 0x1A, 0x21, 0x0B, 0x58, 0x12, 0x23,
	0x2D, 0x24, 0x47, 0x53, 0x19, 0x0C, 0x2A, 0x1A, 0x04, 0x3E, 0x25, 0x2F,
	0x58, 0x4A, 0x0D, 0x2C, 0x14, 0x35, 0x54, 0x57, 0x00, 0x09, 0x19, 0x33,
	0x07, 0x01, 0x03, 0x5B, 0x4E, 0x38, 0x2C, 0x26, 0x43, 0x0C, 0x28, 0x03,
	0x27, 0x55, 0x32, 0x56, 0x44, 0x26, 0x5C, 0x36, 0x02, 0x0D, 0x15, 0x0D,
	0x33, 0x0B, 0x5A, 0x27, 0x47, 0x10, 0x00, 0x3F, 0x69, 0x5E, 0x26, 0x58,
	0x52, 0x0D, 0x5E, 0x03, 0x24, 0x02, 0x23, 0x01, 0x16, 0x0B, 0x2D, 0x6D,
	0x54, 0x16, 0x0D, 0x09, 0x00, 0x22, 0x27, 0x16, 0x02, 0x0D, 0x15, 0x39,
	0x19, 0x2E, 0x0C, 0x02, 0x2E, 0x21, 0x21, 0x13, 0x15, 0x2C, 0x06, 0x0F,
	0x1A, 0x0B, 0x02, 0x0B, 0x39, 0x32, 0x07, 0x56, 0x06, 0x1E, 0x33, 0x06,
	0x35, 0x28, 0x04, 0x33, 0x3E, 0x2B, 0x23, 0x5A, 0x27, 0x20, 0x2B, 0x2B,
	0x5A, 0x14, 0x2E, 0x39, 0x45, 0x1F, 0x00, 0x0A, 0x0C, 0x2C, 0x29, 0x10,
	0x23, 0x4E, 0x1A, 0x0C, 0x24, 0x23, 0x08, 0x5A, 0x28, 0x1B, 0x55, 0x0E,
	0x2D, 0x53, 0x30, 0x1B, 0x26, 0x3B, 0x1C, 0x75, 0x1C, 0x05, 0x3C, 0x07,
	0x05, 0x05, 0x38, 0x23, 0x2E, 0x32, 0x38, 0x2B, 0x04, 0x04, 0x35, 0x29,
	0x34, 0x02, 0x22, 0x0B, 0x59, 0x20, 0x19, 0x18, 0x75, 0x20, 0x0D, 0x1F,
	0x3D, 0x20, 0x2E, 0x59, 0x5C, 0x0E, 0x2D, 0x09, 0x26, 0x09, 0x03, 0x37,
	0x59, 0x24, 0x5D, 0x06, 0x18, 0x5C, 0x22, 0x59, 0x03, 0x23, 0x18, 0x57,
	0x09, 0x02, 0x36, 0x5B, 0x2E, 0x2C, 0x24, 0x2E, 0x5E, 0x06, 0x1C, 0x5C,
	0x3B, 0x54, 0x11, 0x1F, 0x3F, 0x14, 0x1E, 0x0E, 0x36, 0x5F, 0x24, 0x25,
	0x53, 0x07, 0x2F, 0x36, 0x23, 0x27, 0x06, 0x0C, 0x16, 0x08, 0x54, 0x1D,
	0x00, 0x04, 0x23, 0x0A, 0x0A, 0x40, 0x12, 0x3F, 0x07, 0x0F, 0x44, 0x15,
	0x03, 0x02, 0x21, 0x04, 0x2D, 0x2F, 0x2E, 0x19, 0x40, 0x28, 0x09, 0x0D,
	0x1D, 0x25, 0x1A, 0x28, 0x36, 0x0B, 0x40, 0x6D, 0x3E, 0x13, 0x5B, 0x58,
	0x1A, 0x15, 0x34, 0x1D, 0x3C, 0x35, 0x00, 0x4A, 0x27, 0x20, 0x71, 0x3A,
	0x18, 0x0A, 0x5A, 0x37, 0x18, 0x28, 0x37, 0x27, 0x7B, 0x24, 0x35, 0x20,
	0x20, 0x05, 0x16, 0x35, 0x08, 0x5A, 0x2D, 0x04, 0x04, 0x59, 0x1B, 0x00,
	0x21, 0x57, 0x14, 0x26, 0x75, 0x1C, 0x55, 0x3A, 0x1F, 0x05, 0x06, 0x26,
	0x37, 0x58, 0x0C, 0x0E, 0x0E, 0x0D, 0x1A, 0x29, 0x24, 0x08, 0x1C, 0x1A,
	0x00, 0x54, 0x0A, 0x37, 0x20, 0x21, 0x2B, 0x10, 0x1F, 0x5A, 0x24, 0x5C,
	0x2D, 0x22, 0x1F, 0x3B, 0x0F, 0x03, 0x2C, 0x12, 0x7B, 0x09, 0x2A, 0x1C,
	0x2D, 0x73, 0x5C, 0x37, 0x1C, 0x2D, 0x33, 0x54, 0x4E, 0x25, 0x1A, 0x04,
	0x47, 0x11, 0x3B, 0x18, 0x1A, 0x1E, 0x24, 0x01, 0x20, 0x72, 0x5E, 0x0A,
	0x0D, 0x1C, 0x0C, 0x3B, 0x2B, 0x02, 0x0F, 0x0A, 0x35, 0x04, 0x1A, 0x20,
	0x0F, 0x19, 0x0B, 0x24, 0x5D, 0x29, 0x5C, 0x18, 0x03, 0x07, 0x30, 0x2A,
	0x32, 0x06, 0x3A, 0x2F, 0x1D, 0x34, 0x27, 0x3C, 0x18, 0x34, 0x2E, 0x23,
	0x03, 0x00, 0x21, 0x55, 0x21, 0x52, 0x24, 0x2A, 0x32, 0x26, 0x25, 0x2D,
	0x18, 0x23, 0x3A, 0x21, 0x71, 0x43, 0x32, 0x5D, 0x22, 0x17, 0x22, 0x07,
	0x18, 0x33, 0x08, 0x00, 0x2C, 0x2C, 0x3E, 0x76, 0x0B, 0x38, 0x3B, 0x3B,
	0x34, 0x1E, 0x33, 0x3D, 0x23, 0x09, 0x15, 0x1B, 0x2B, 0x1D, 0x00, 0x24,
	0x2C, 0x56, 0x3E, 0x74, 0x0A, 0x51, 0x41, 0x44, 0x73, 0x27, 0x55, 0x00,
	0x0E, 0x07, 0x25, 0x03, 0x57, 0x28, 0x3A, 0x0A, 0x0F, 0x0F, 0x3F, 0x33,
	0x5A, 0x27, 0x0A, 0x44, 0x31, 0x34, 0x13, 0x24, 0x2D, 0x3B, 0x19, 0x0B,
	0x04, 0x19, 0x75, 0x2D, 0x2F, 0x34, 0x12, 0x77, 0x3E, 0x33, 0x3E, 0x44,
	0x0F, 0x07, 0x57, 0x5E, 0x3C, 0x21, 0x28, 0x0F, 0x2F, 0x2A, 0x14, 0x34,
	0x34, 0x3E, 0x0F, 0x21, 0x19, 0x05, 0x06, 0x53, 0x21, 0x47, 0x4E, 0x36,
	0x29, 0x21, 0x21, 0x13, 0x0A, 0x28, 0x74, 0x26, 0x17, 0x04, 0x13, 0x0C,
	0x05, 0x2E, 0x37, 0x3B, 0x14, 0x16, 0x33, 0x0F, 0x53, 0x72, 0x5D, 0x20,
	0x2B, 0x44, 0x69, 0x58, 0x0A, 0x2B, 0x5B, 0x23, 0x5B, 0x51, 0x1F, 0x53,
	0x0D, 0x2A, 0x19, 0x09, 0x06, 0x18, 0x3B, 0x2D, 0x26, 0x0E, 0x77, 0x00,
	0x51, 0x37, 0x1B, 0x05, 0x5F, 0x39, 0x0F, 0x18, 0x18, 0x0A, 0x36, 0x28,
	0x24, 0x30, 0x27, 0x15, 0x2C, 0x21, 0x0E, 0x1E, 0x09, 0x18, 0x3D, 0x70,
	0x06, 0x37, 0x20, 0x44, 0x37, 0x25, 0x15, 0x39, 0x20, 0x75, 0x5E, 0x15,
	0x37, 0x06, 0x36, 0x35, 0x35, 0x0F, 0x02, 0x12, 0x21, 0x14, 0x2B, 0x1F,
	0x3B, 0x34, 0x2D, 0x22, 0x11, 0x32, 0x03, 0x1B, 0x5A, 0x08, 0x09, 0x58,
	0x51, 0x0B, 0x32, 0x38, 0x3F, 0x37, 0x39, 0x38, 0x16, 0x04, 0x25, 0x37,
	0x3F, 0x01, 0x3C, 0x1B, 0x0F, 0x5E, 0x08, 0x59, 0x11, 0x29, 0x32, 0x74,
	0x08, 0x10, 0x03, 0x5B, 0x6D, 0x5A, 0x02, 0x17, 0x1D, 0x18, 0x22, 0x07,
	0x3D, 0x3E, 0x2E, 0x19, 0x00, 0x02, 0x0D, 0x0B, 0x3D, 0x27, 0x0C, 0x27,
	0x34, 0x14, 0x51, 0x17, 0x02, 0x05, 0x06, 0x12, 0x1A, 0x2F, 0x2F, 0x27,
	0x35, 0x0F, 0x24, 0x3A, 0x3B, 0x08, 0x5E, 0x2E, 0x10, 0x3A, 0x56, 0x3B,
	0x3D, 0x24, 0x26, 0x10, 0x45, 0x06, 0x2B, 0x5C, 0x55, 0x5C, 0x32, 0x75,
	0x22, 0x08, 0x1C, 0x33, 0x28, 0x1A, 0x12, 0x09, 0x58, 0x31, 0x27, 0x31,
	0x3E, 0x08, 0x12, 0x5B, 0x07, 0x0F, 0x09, 0x71, 0x09, 0x54, 0x3A, 0x40,
	0x16, 0x01, 0x2F, 0x1D, 0x28, 0x7A, 0x5E, 0x09, 0x2D, 0x3D, 0x03, 0x19,
	0x25, 0x02, 0x0D, 0x14, 0x07, 0x0A, 0x34, 0x59, 0x18, 0x00, 0x36, 0x56,
	0x03, 0x13, 0x22, 0x4E, 0x00, 0x23, 0x07, 0x38, 0x58, 0x2F, 0x59, 0x18,
	0x55, 0x03, 0x00, 0x2A, 0x32, 0x2E, 0x4E, 0x1E, 0x04, 0x27, 0x0D, 0x0D,
	0x26, 0x1A, 0x2C, 0x54, 0x30, 0x2C, 0x5B, 0x74, 0x06, 0x36, 0x17, 0x06,
	0x2F, 0x58, 0x57, 0x0D, 0x21, 0x30, 0x54, 0x53, 0x5B, 0x0A, 0x7B, 0x27,
	0x18, 0x5E, 0x5B, 0x2C, 0x34, 0x53, 0x41, 0x59, 0x08, 0x0E, 0x1B, 0x41,
	0x0D, 0x72, 0x19, 0x0D, 0x1F, 0x3F, 0x15, 0x2B, 0x39, 0x02, 0x09, 0x13,
	0x2B, 0x0F, 0x0A, 0x1C, 0x14, 0x19, 0x24, 0x56, 0x58, 0x0E, 0x2E, 0x51,
	0x0F, 0x3D, 0x3B, 0x55, 0x12, 0x0C, 0x5E, 0x23, 0x20, 0x22, 0x21, 0x40,
	0x32, 0x2A, 0x03, 0x58, 0x13, 0x06, 0x1B, 0x00, 0x20, 0x5F, 0x2D, 0x0F,
	0x39, 0x59, 0x29, 0x18, 0x36, 0x23, 0x39, 0x24, 0x74, 0x22, 0x04, 0x04,
	0x38, 0x2D, 0x01, 0x29, 0x45, 0x32, 0x18, 0x0D, 0x0A, 0x58, 0x24, 0x05,
	0x59, 0x2D, 0x28, 0x33, 0x7B, 0x36, 0x0B, 0x38, 0x3D, 0x73, 0x43, 0x34,
	0x0C, 0x1E, 0x2C, 0x03, 0x3B, 0x58, 0x5A, 0x11, 0x0D, 0x11, 0x03, 0x5F,
	0x13, 0x2B, 0x2B, 0x29, 0x5B, 0x12, 0x43, 0x39, 0x58, 0x2C, 0x20, 0x2F,
	0x17, 0x1D, 0x19, 0x2F, 0x38, 0x29, 0x0D, 0x07, 0x3B, 0x1B, 0x27, 0x16,
	0x23, 0x12, 0x2F, 0x2A, 0x18, 0x01, 0x29, 0x5D, 0x55, 0x36, 0x21, 0x72,
	0x1B, 0x09, 0x37, 0x3B, 0x2F, 0x16, 0x50, 0x22, 0x40, 0x0D, 0x01, 0x58,
	0x02, 0x33, 0x33, 0x06, 0x33, 0x1A, 0x53, 0x37, 0x18, 0x3B, 0x41, 0x5E,
	0x26, 0x34, 0x2C, 0x05, 0x19, 0x07, 0x58, 0x17, 0x22, 0x0E, 0x2B, 0x04,
	0x39, 0x5F, 0x0A, 0x20, 0x34, 0x50, 0x3A, 0x0E, 0x13, 0x3A, 0x53, 0x26,
	0x5E, 0x2F, 0x3C, 0x16, 0x5C, 0x2A, 0x37, 0x0F, 0x56, 0x23, 0x28, 0x34,
	0x1D, 0x57, 0x0B, 0x13, 0x15, 0x04, 0x37, 0x0F, 0x5F, 0x32, 0x43, 0x15,
	0x26, 0x38, 0x28, 0x1E, 0x30, 0x3B, 0x33, 0x0A, 0x24, 0x36, 0x1F, 0x5A,
	0x08, 0x02, 0x33, 0x45, 0x1F, 0x0C, 0x5A, 0x52, 0x34, 0x21, 0x71, 0x2B,
	0x24, 0x38, 0x08, 0x73, 0x5A, 0x07, 0x26, 0x19, 0x1A, 0x04, 0x37, 0x29,
	0x09, 0x15, 0x26, 0x2E, 0x02, 0x5E, 0x2C, 0x03, 0x23, 0x04, 0x08, 0x17,
	0x2E, 0x55, 0x1A, 0x59, 0x07, 0x39, 0x34, 0x18, 0x0A, 0x15, 0x04, 0x14,
	0x18, 0x0C, 0x34, 0x16, 0x0A, 0x0D, 0x1C, 0x10, 0x35, 0x59, 0x26, 0x22,
	0x09, 0x00, 0x51, 0x22, 0x18, 0x6D, 0x0D, 0x2B, 0x17, 0x11, 0x2D, 0x3A,
	0x0D, 0x0B, 0x08, 0x74, 0x5E, 0x58, 0x36, 0x09, 0x71, 0x38, 0x1B, 0x27,
	0x02, 0x2E, 0x3A, 0x32, 0x27, 0x0C, 0x17, 0x5F, 0x37, 0x20, 0x31, 0x33,
	0x0F, 0x25, 0x01, 0x07, 0x37, 0x39, 0x19, 0x57, 0x20, 0x37, 0x14, 0x0A,
	0x36, 0x04, 0x13, 0x26, 0x32, 0x2C, 0x3F, 0x2D, 0x0D, 0x06, 0x18, 0x1B,
	0x3A, 0x16, 0x38, 0x57, 0x2F, 0x11, 0x1A, 0x20, 0x20, 0x3C, 0x13, 0x1E,
	0x59, 0x3F, 0x21, 0x74, 0x34, 0x04, 0x38, 0x12, 0x2C, 0x03, 0x4A, 0x14,
	0x31, 0x7B, 0x23, 0x27, 0x2F, 0x07, 0x12, 0x03, 0x20, 0x0D, 0x58, 0x0F,
	0x3D, 0x0B, 0x1A, 0x24, 0x04, 0x16, 0x08, 0x01, 0x01, 0x7B, 0x18, 0x16,
	0x1D, 0x22, 0x75, 0x2B, 0x09, 0x14, 0x04, 0x2F, 0x5C, 0x57, 0x59, 0x5A,
	0x72, 0x04, 0x35, 0x2A, 0x1F, 0x28, 0x04, 0x33, 0x2C, 0x04, 0x12, 0x5A,
	0x2D, 0x03, 0x58, 0x25, 0x39, 0x4E, 0x41, 0x02, 0x06, 0x2D, 0x33, 0x1C,
	0x04, 0x29, 0x3B, 0x57, 0x19, 0x52, 0x33, 0x1A, 0x51, 0x1A, 0x22, 0x30,
	0x1E, 0x00, 0x1E, 0x01, 0x07, 0x54, 0x32, 0x57, 0x05, 0x05, 0x0F, 0x20,
	0x45, 0x1B, 0x15, 0x24, 0x30, 0x16, 0x38, 0x1A, 0x27, 0x16, 0x5C, 0x0F,
	0x23, 0x00, 0x12, 0x00, 0x2E, 0x7B, 0x5C, 0x2E, 0x41, 0x3B, 0x0F, 0x3C,
	0x39, 0x21, 0x19, 0x03, 0x0D, 0x2F, 0x3C, 0x04, 0x36, 0x5C, 0x0E, 0x06,
	0x23, 0x7A, 0x15, 0x10, 0x19, 0x06, 0x15, 0x2A, 0x0A, 0x3F, 0x13, 0x3A,
	0x3A, 0x30, 0x3E, 0x3B, 0x12, 0x25, 0x1B, 0x5C, 0x0F, 0x1A, 0x02, 0x52,
	0x39, 0x03, 0x09, 0x55, 0x34, 0x21, 0x2E, 0x01, 0x22, 0x37, 0x05, 0x1A,
	0x34, 0x58, 0x38, 0x5E, 0x31, 0x05, 0x3D, 0x4A, 0x1D, 0x18, 0x33, 0x5D,
	0x26, 0x3D, 0x05, 0x37, 0x3B, 0x56, 0x2A, 0x5E, 0x0F, 0x2F, 0x38, 0x20,
	0x3E, 0x04, 0x18, 0x04, 0x21, 0x07, 0x35, 0x5C, 0x36, 0x20, 0x2D, 0x37,
	0x1E, 0x08, 0x34, 0x39, 0x3B, 0x47, 0x2F, 0x0D, 0x0E, 0x30, 0x15, 0x39,
	0x24, 0x07, 0x38, 0x5A, 0x4E, 0x5A, 0x5A, 0x2A, 0x1D, 0x19, 0x5B, 0x3C,
	0x69, 0x3B, 0x09, 0x34, 0x0A, 0x31, 0x3E, 0x1B, 0x5D, 0x05, 0x35, 0x3A,
	0x23, 0x1C, 0x31, 0x06, 0x00, 0x22, 0x0B, 0x0D, 0x11, 0x02, 0x58, 0x0A,
	0x27, 0x1A, 0x1D, 0x0E, 0x03, 0x3A, 0x36, 0x0A, 0x32, 0x59, 0x5A, 0x20,
	0x24, 0x34, 0x38, 0x00, 0x2E, 0x04, 0x1B, 0x3B, 0x0A, 0x73, 0x01, 0x3B,
	0x2C, 0x24, 0x24, 0x27, 0x27, 0x39, 0x5A, 0x03, 0x04, 0x04, 0x34, 0x21,
	0x14, 0x03, 0x02, 0x16, 0x0F, 0x76, 0x47, 0x37, 0x21, 0x01, 0x2B, 0x0A,
	0x00, 0x25, 0x3E, 0x2F, 0x14, 0x4E, 0x1D, 0x2C, 0x09, 0x15, 0x51, 0x0F,
	0x2F, 0x15, 0x59, 0x56, 0x18, 0x0F, 0x17, 0x04, 0x34, 0x22, 0x2E, 0x7B,
	0x29, 0x59, 0x26, 0x06, 0x24, 0x04, 0x59, 0x1D, 0x08, 0x33, 0x16, 0x25,
	0x34, 0x29, 0x2A, 0x0F, 0x51, 0x0F, 0x5E, 0x15, 0x3A, 0x58, 0x24, 0x52,
	0x2F, 0x35, 0x57, 0x1C, 0x5F, 0x05, 0x3D, 0x10, 0x3B, 0x3B, 0x75, 0x0E,
	0x0A, 0x28, 0x5D, 0x11, 0x5C, 0x51, 0x1B, 0x0C, 0x11, 0x39, 0x4E, 0x38,
	0x1B, 0x2A, 0x1A, 0x52, 0x1D, 0x59, 0x0E, 0x0F, 0x18, 0x38, 0x5B, 0x2C,
	0x1D, 0x55, 0x23, 0x06, 0x05, 0x3C, 0x51, 0x2C, 0x38, 0x0E, 0x5F, 0x36,
	0x3A, 0x0F, 0x11, 0x0E, 0x02, 0x14, 0x31, 0x76, 0x07, 0x37, 0x25, 0x33,
	0x21, 0x22, 0x2C, 0x0A, 0x1C, 0x12, 0x05, 0x25, 0x0B, 0x0C, 0x77, 0x23,
	0x09, 0x02, 0x08, 0x7B, 0x1C, 0x0C, 0x03, 0x38, 0x3A, 0x01, 0x2F, 0x57,
	0x59, 0x12, 0x0B, 0x3B, 0x5B, 0x0C, 0x18, 0x5D, 0x35, 0x1A, 0x0A, 0x2B,
	0x2F, 0x0F, 0x03, 0x18, 0x0C, 0x29, 0x34, 0x23, 0x19, 0x77, 0x2A, 0x0B,
	0x02, 0x0F, 0x0C, 0x39, 0x32, 0x3B, 0x2D, 0x73, 0x5E, 0x19, 0x5E, 0x5E,
	0x27, 0x1E, 0x34, 0x0A, 0x1E, 0x2E, 0x05, 0x0B, 0x14, 0x0F, 0x69, 0x34,
	0x2B, 0x1A, 0x0C, 0x70, 0x5F, 0x16, 0x5C, 0x1D, 0x34, 0x21, 0x07, 0x2A,
	0x0F, 0x2C, 0x23, 0x0A, 0x2D, 0x18, 0x30, 0x0D, 0x57, 0x1A, 0x24, 0x74,
	0x1A, 0x33, 0x5A, 0x5E, 0x20, 0x2A, 0x02, 0x01, 0x19, 0x76, 0x18, 0x4E,
	0x59, 0x0A, 0x7B, 0x00, 0x24, 0x03, 0x1F, 0x2C, 0x3B, 0x22, 0x0B, 0x03,
	0x33, 0x0D, 0x16, 0x0C, 0x27, 0x72, 0x02, 0x28, 0x26, 0x32, 0x13, 0x28,
	0x20, 0x59, 0x3D, 0x23, 0x2A, 0x2E, 0x26, 0x25, 0x08, 0x09, 0x57, 0x07,
	0x24, 0x20, 0x29, 0x0D, 0x25, 0x07, 0x1A, 0x54, 0x30, 0x0A, 0x09, 0x18,
	0x24, 0x34, 0x17, 0x0F, 0x07, 0x00, 0x57, 0x3D, 0x20, 0x01, 0x14, 0x36,
	0x2D, 0x52, 0x15, 0x20, 0x05, 0x3B, 0x44, 0x2A, 0x54, 0x2F, 0x38, 0x1A,
	0x6D, 0x0E, 0x0F, 0x39, 0x01, 0x0D, 0x3D, 0x05, 0x0B, 0x1E, 0x34, 0x5B,
	0x17, 0x28, 0x1B, 0x04, 0x0A, 0x35, 0x58, 0x31, 0x15, 0x03, 0x19, 0x08,
	0x58, 0x0D, 0x5B, 0x53, 0x24, 0x11, 0x6D, 0x5A, 0x10, 0x3E, 0x3F, 0x03,
	0x3A, 0x33, 0x1F, 0x3A, 0x18, 0x0B, 0x2A, 0x05, 0x1D, 0x2C, 0x19, 0x50,
	0x36, 0x0F, 0x00, 0x36, 0x03, 0x21, 0x5A, 0x2A, 0x5A, 0x0A, 0x22, 0x08,
	0x29, 0x0E, 0x36, 0x58, 0x3D, 0x16, 0x00, 0x30, 0x06, 0x08, 0x04, 0x2B,
	0x11, 0x0F, 0x11, 0x17, 0x00, 0x0A, 0x58, 0x5D, 0x11, 0x06, 0x10, 0x0F,
	0x24, 0x30, 0x08, 0x03, 0x59, 0x3F, 0x15, 0x18, 0x0A, 0x09, 0x53, 0x04,
	0x0E, 0x55, 0x01, 0x53, 0x35, 0x02, 0x55, 0x0B, 0x1B, 0x34, 0x3E, 0x29,
	0x28, 0x3D, 0x21, 0x1D, 0x39, 0x2B, 0x23, 0x74, 0x25, 0x2E, 0x1A, 0x31,
	0x75, 0x3F, 0x28, 0x5E, 0x59, 0x13, 0x0D, 0x2B, 0x37, 0x3D, 0x09, 0x19,
	0x33, 0x24, 0x1C, 0x00, 0x3A, 0x58, 0x3C, 0x1E, 0x09, 0x0F, 0x04, 0x1C,
	0x44, 0x0F, 0x19, 0x39, 0x09, 0x19, 0x08, 0x0D, 0x24, 0x00, 0x3B, 0x06,
	0x47, 0x24, 0x20, 0x07, 0x29, 0x1B, 0x0C, 0x04, 0x19, 0x00, 0x3E, 0x17,
	0x5B, 0x23, 0x0E, 0x1D, 0x0A, 0x14, 0x26, 0x1A, 0x1D, 0x15, 0x3B, 0x5A,
	0x29, 0x5E, 0x0B, 0x2D, 0x0D, 0x33, 0x47, 0x0F, 0x34, 0x31, 0x14, 0x24,
	0x24, 0x59, 0x1A, 0x0E, 0x3E, 0x31, 0x59, 0x00, 0x11, 0x09, 0x31, 0x3E,
	0x0F, 0x0A, 0x1C, 0x1B, 0x3F, 0x02, 0x77, 0x24, 0x08, 0x0B, 0x02, 0x70,
	0x09, 0x3B, 0x24, 0x59, 0x0D, 0x14, 0x59, 0x20, 0x5A, 0x72, 0x04, 0x29,
	0x2C, 0x5D, 0x2C, 0x06, 0x0C, 0x5F, 0x00, 0x7B, 0x5F, 0x2F, 0x16, 0x3E,
	0x05, 0x3D, 0x50, 0x24, 0x13, 0x25, 0x19, 0x58, 0x1C, 0x21, 0x08, 0x27,
	0x04, 0x3E, 0x2C, 0x1A, 0x3C, 0x23, 0x1D, 0x1F, 0x34, 0x0A, 0x3B, 0x59,
	0x58, 0x31, 0x1F, 0x57, 0x3D, 0x52, 0x09, 0x29, 0x2C, 0x1B, 0x19, 0x38,
	0x01, 0x13, 0x04, 0x0C, 0x2F, 0x5A, 0x53, 0x37, 0x38, 0x27, 0x43, 0x2F,
	0x3A, 0x0A, 0x29, 0x5A, 0x2F, 0x56, 0x1F, 0x36, 0x28, 0x35, 0x25, 0x26,
	0x33, 0x29, 0x04, 0x5E, 0x5F, 0x77, 0x26, 0x58, 0x08, 0x1C, 0x12, 0x2A,
	0x00, 0x23, 0x2F, 0x32, 0x5C, 0x24, 0x0F, 0x19, 0x0C, 0x1A, 0x13, 0x58,
	0x2A, 0x30, 0x23, 0x34, 0x1C, 0x2D, 0x1B, 0x1F, 0x18, 0x24, 0x1C, 0x33,
	0x3B, 0x00, 0x5E, 0x0D, 0x0C, 0x5A, 0x11, 0x1E, 0x25, 0x33, 0x27, 0x00,
	0x26, 0x3D, 0x16, 0x2F, 0x0D, 0x39, 0x31, 0x2D, 0x5D, 0x59, 0x05, 0x2A,
	0x15, 0x5C, 0x53, 0x2A, 0x24, 0x01, 0x14, 0x07, 0x0F, 0x0E, 0x31, 0x28,
	0x36, 0x2C, 0x1D, 0x0B, 0x15, 0x57, 0x1E, 0x22, 0x26, 0x09, 0x33, 0x07,
	0x26, 0x30, 0x39, 0x39, 0x20, 0x18, 0x33, 0x04, 0x4A, 0x0D, 0x13, 0x15,
	0x43, 0x50, 0x25, 0x01, 0x18, 0x1D, 0x39, 0x0D, 0x1A, 0x17, 0x08, 0x57,
	0x07, 0x04, 0x15, 0x5B, 0x22, 0x34, 0x1E, 0x2F, 0x3B, 0x15, 0x5E, 0x1F,
	0x07, 0x3F, 0x0D, 0x5C, 0x52, 0x25, 0x58, 0x55, 0x2D, 0x25, 0x00, 0x39,
	0x18, 0x59, 0x29, 0x08, 0x5D, 0x11, 0x07, 0x19, 0x75, 0x5F, 0x06, 0x5A,
	0x3C, 0x00, 0x3B, 0x15, 0x28, 0x11, 0x75, 0x08, 0x39, 0x1A, 0x00, 0x1A,
	0x39, 0x07, 0x56, 0x0A, 0x17, 0x2B, 0x38, 0x1A, 0x44, 0x75, 0x1D, 0x11,
	0x5D, 0x0E, 0x06, 0x5C, 0x3B, 0x56, 0x33, 0x05, 0x09, 0x15, 0x09, 0x1E,
	0x0F, 0x00, 0x15, 0x0A, 0x07, 0x0F, 0x58, 0x12, 0x5C, 0x0C, 0x32, 0x0D,
	0x37, 0x1A, 0x0D, 0x70, 0x0B, 0x31, 0x22, 0x1A, 0x72, 0x1A, 0x0D, 0x28,
	0x09, 0x75, 0x34, 0x33, 0x59, 0x12, 0x76, 0x01, 0x2F, 0x17, 0x33, 0x01,
	0x36, 0x20, 0x5B, 0x33, 0x1A, 0x24, 0x59, 0x27, 0x0F, 0x16, 0x1A, 0x0A,
	0x58, 0x2D, 0x24, 0x0E, 0x13, 0x39, 0x0A, 0x15, 0x5A, 0x00, 0x5C, 0x05,
	0x76, 0x08, 0x09, 0x05, 0x1D, 0x05, 0x3B, 0x27, 0x17, 0x03, 0x12, 0x06,
	0x03, 0x1D, 0x5E, 0x31, 0x36, 0x16, 0x27, 0x58, 0x73, 0x47, 0x28, 0x1E,
	0x02, 0x14, 0x22, 0x4E, 0x06, 0x07, 0x16, 0x15, 0x13, 0x3A, 0x5C, 0x27,
	0x19, 0x02, 0x01, 0x24, 0x14, 0x2A, 0x16, 0x01, 0x1B, 0x21, 0x29, 0x12,
	0x0F, 0x44, 0x74, 0x35, 0x2A, 0x3B, 0x5A, 0x77, 0x23, 0x57, 0x58, 0x03,
	0x32, 0x3F, 0x28, 0x1A, 0x11, 0x05, 0x04, 0x04, 0x29, 0x27, 0x7B, 0x1B,
	0x05, 0x3D, 0x0A, 0x73, 0x47, 0x33, 0x06, 0x21, 0x24, 0x04, 0x16, 0x1E,
	0x1F, 0x1A, 0x26, 0x28, 0x1A, 0x5A, 0x29, 0x5E, 0x0D, 0x5F, 0x19, 0x27,
	0x27, 0x2B, 0x0F, 0x33, 0x23, 0x54, 0x58, 0x17, 0x3F, 0x16, 0x26, 0x17,
	0x1A, 0x32, 0x32, 0x28, 0x04, 0x1B, 0x5F, 0x09, 0x2D, 0x09, 0x3B, 0x5A,
	0x31, 0x08, 0x2E, 0x1B, 0x3C, 0x2C, 0x15, 0x19, 0x5C, 0x3E, 0x28, 0x5C,
	0x29, 0x21, 0x5A, 0x74, 0x06, 0x07, 0x1F, 0x02, 0x73, 0x0D, 0x24, 0x3C,
	0x20, 0x1B, 0x2F, 0x09, 0x1D, 0x21, 0x17, 0x23, 0x4E, 0x38, 0x31, 0x0B,
	0x5E, 0x12, 0x09, 0x2C, 0x00, 0x29, 0x04, 0x37, 0x33, 0x05, 0x0E, 0x2E,
	0x1D, 0x09, 0x27, 0x36, 0x3B, 0x2B, 0x58, 0x09, 0x36, 0x52, 0x3E, 0x2C,
	0x1B, 0x19, 0x03, 0x29, 0x22, 0x08, 0x3A, 0x2F, 0x16, 0x21, 0x74, 0x1F,
	0x26, 0x38, 0x08, 0x72, 0x0D, 0x12, 0x09, 0x20, 0x0E, 0x27, 0x09, 0x2C,
	0x09, 0x1A, 0x36, 0x12, 0x56, 0x3F, 0x3B, 0x0B, 0x15, 0x5C, 0x1C, 0x77,
	0x1D, 0x4A, 0x41, 0x31, 0x08, 0x06, 0x29, 0x0A, 0x01, 0x28, 0x3B, 0x0D,
	0x21, 0x02, 0x11, 0x0E, 0x00, 0x57, 0x25, 0x09, 0x5A, 0x4E, 0x1A, 0x2C,
	0x3B, 0x0D, 0x18, 0x1E, 0x5D, 0x2A, 0x15, 0x0A, 0x5B, 0x05, 0x00, 0x20,
	0x53, 0x0A, 0x5E, 0x0D, 0x34, 0x19, 0x59, 0x0C, 0x15, 0x25, 0x37, 0x5C,
	0x04, 0x70, 0x1A, 0x27, 0x5E, 0x04, 0x00, 0x47, 0x13, 0x41, 0x04, 0x38,
	0x1F, 0x15, 0x21, 0x1B, 0x28, 0x3F, 0x53, 0x58, 0x2C, 0x04, 0x07, 0x57,
	0x57, 0x28, 0x27, 0x38, 0x2C, 0x59, 0x59, 0x25, 0x1F, 0x39, 0x02, 0x40,
	0x2D, 0x34, 0x2E, 0x23, 0x2F, 0x70, 0x15, 0x34, 0x41, 0x04, 0x18, 0x23,
	0x52, 0x27, 0x18, 0x20, 0x0F, 0x0A, 0x5F, 0x3C, 0x6D, 0x3A, 0x18, 0x1D,
	0x53, 0x38, 0x23, 0x53, 0x5B, 0x53, 0x3B, 0x01, 0x26, 0x5A, 0x0C, 0x70,
	0x15, 0x0C, 0x2D, 0x05, 0x15, 0x34, 0x23, 0x3C, 0x24, 0x17, 0x00, 0x26,
	0x20, 0x39, 0x37, 0x5B, 0x52, 0x3C, 0x3F, 0x33, 0x5D, 0x16, 0x0C, 0x2F,
	0x31, 0x01, 0x06, 0x3C, 0x1D, 0x69, 0x24, 0x4A, 0x1D, 0x27, 0x15, 0x3F,
	0x37, 0x2D, 0x13, 0x0C, 0x3E, 0x02, 0x34, 0x07, 0x26, 0x24, 0x32, 0x1B,
	0x2C, 0x16, 0x47, 0x50, 0x04, 0x0A, 0x1B, 0x54, 0x0E, 0x3F, 0x19, 0x01,
	0x3B, 0x57, 0x08, 0x31, 0x18, 0x1A, 0x2F, 0x0F, 0x05, 0x10, 0x09, 0x27,
	0x5F, 0x09, 0x75, 0x21, 0x2D, 0x1E, 0x2E, 0x76, 0x26, 0x2D, 0x5A, 0x29,
	0x14, 0x1D, 0x51, 0x00, 0x23, 0x2A, 0x3A, 0x29, 0x06, 0x03, 0x3A, 0x5B,
	0x32, 0x3F, 0x53, 0x29, 0x5B, 0x0F, 0x41, 0x18, 0x13, 0x1B, 0x4A, 0x3A,
	0x21, 0x34, 0x27, 0x56, 0x08, 0x3E, 0x34, 0x02, 0x27, 0x5F, 0x0E, 0x0F,
	0x16, 0x03, 0x0B, 0x29, 0x08, 0x07, 0x26, 0x1A, 0x3F, 0x0D, 0x15, 0x13,
	0x01, 0x3B, 0x7A, 0x5C, 0x36, 0x08, 0x44, 0x71, 0x5C, 0x19, 0x57, 0x20,
	0x75, 0x35, 0x08, 0x3A, 0x06, 0x37, 0x34, 0x02, 0x1E, 0x1D, 0x08, 0x0E,
	0x57, 0x28, 0x26, 0x2C, 0x2B, 0x00, 0x57, 0x03, 0x30, 0x24, 0x53, 0x58,
	0x03, 0x15, 0x38, 0x39, 0x56, 0x3C, 0x03, 0x5D, 0x55, 0x02, 0x04, 0x10,
	0x1D, 0x10, 0x2C, 0x1C, 0x0F, 0x1F, 0x2F, 0x5F, 0x3C, 0x29, 0x54, 0x28,
	0x5A, 0x40, 0x17, 0x07, 0x11, 0x59, 0x1A, 0x17, 0x09, 0x35, 0x3A, 0x58,
	0x76, 0x16, 0x14, 0x1F, 0x21, 0x2B, 0x20, 0x4E, 0x06, 0x3B, 0x72, 0x27,
	0x13, 0x34, 0x19, 0x11, 0x3B, 0x2A, 0x06, 0x20, 0x34, 0x5B, 0x23, 0x39,
	0x26, 0x7B, 0x1F, 0x29, 0x08, 0x26, 0x71, 0x39, 0x19, 0x34, 0x5B, 0x24,
	0x3B, 0x02, 0x0B, 0x58, 0x29, 0x5C, 0x50, 0x22, 0x2D, 0x31, 0x54, 0x37,
	0x3D, 0x07, 0x07, 0x0D, 0x55, 0x04, 0x33, 0x70, 0x14, 0x04, 0x05, 0x22,
	0x2C, 0x2E, 0x56, 0x5D, 0x5E, 0x2E, 0x2E, 0x1B, 0x58, 0x5E, 0x2B, 0x5E,
	0x30, 0x1F, 0x3D, 0x7A, 0x36, 0x29, 0x3D, 0x29, 0x12, 0x1E, 0x07, 0x21,
	0x23, 0x27, 0x24, 0x30, 0x2F, 0x22, 0x26, 0x3A, 0x00, 0x3F, 0x0A, 0x09,
	0x3A, 0x31, 0x04, 0x25, 0x23, 0x2D, 0x59, 0x41, 0x1F, 0x21, 0x38, 0x2E,
	0x1B, 0x33, 0x2D, 0x1B, 0x57, 0x1A, 0x22, 0x20, 0x25, 0x53, 0x5A, 0x33,
	0x3B, 0x43, 0x20, 0x58, 0x0A, 0x30, 0x22, 0x32, 0x1B, 0x5B, 0x74, 0x2A,
	0x00, 0x5E, 0x59, 0x72, 0x24, 0x22, 0x37, 0x13, 0x0B, 0x03, 0x18, 0x5B,
	0x38, 0x27, 0x1E, 0x12, 0x03, 0x19, 0x01, 0x5C, 0x0C, 0x41, 0x53, 0x13,
	0x22, 0x1B, 0x0F, 0x2C, 0x18, 0x26, 0x54, 0x5D, 0x32, 0x21, 0x26, 0x0A,
	0x06, 0x5E, 0x75, 0x1F, 0x54, 0x2C, 0x40, 0x38, 0x34, 0x3B, 0x06, 0x40,
	0x3B, 0x58, 0x30, 0x04, 0x52, 0x27, 0x0E, 0x50, 0x3F, 0x3A, 0x24, 0x01,
	0x50, 0x5E, 0x1A, 0x29, 0x2A, 0x36, 0x36, 0x59, 0x2F, 0x03, 0x59, 0x3A,
	0x03, 0x37, 0x2D, 0x33, 0x3D, 0x29, 0x73, 0x3F, 0x33, 0x0B, 0x18, 0x09,
	0x36, 0x0C, 0x5F, 0x2D, 0x18, 0x16, 0x10, 0x5E, 0x12, 0x18, 0x2D, 0x53,
	0x27, 0x3F, 0x08, 0x35, 0x26, 0x3C, 0x52, 0x32, 0x16, 0x35, 0x41, 0x0C,
	0x2F, 0x26, 0x17, 0x17, 0x29, 0x74, 0x0B, 0x1B, 0x5E, 0x5C, 0x13, 0x34,
	0x51, 0x3A, 0x39, 0x0B, 0x0E, 0x19, 0x24, 0x26, 0x2F, 0x3F, 0x0E, 0x26,
	0x26, 0x74, 0x05, 0x50, 0x58, 0x5D, 0x04, 0x0D, 0x54, 0x17, 0x07, 0x0C,
	0x2E, 0x4A, 0x27, 0x5E, 0x25, 0x04, 0x58, 0x25, 0x5E, 0x13, 0x25, 0x52,
	0x45, 0x18, 0x38, 0x2F, 0x31, 0x18, 0x1D, 0x16, 0x2A, 0x35, 0x20, 0x0F,
	0x10, 0x27, 0x26, 0x36, 0x33, 0x7A, 0x5B, 0x2E, 0x1F, 0x25, 0x0E, 0x24,
	0x3B, 0x3E, 0x32, 0x73, 0x1D, 0x53, 0x3F, 0x1A, 0x21, 0x5B, 0x05, 0x5F,
	0x44, 0x14, 0x27, 0x03, 0x39, 0x1A, 0x08, 0x16, 0x08, 0x14, 0x1E, 0x0F,
	0x3D, 0x0B, 0x37, 0x13, 0x69, 0x3D, 0x31, 0x16, 0x5A, 0x2D, 0x14, 0x12,
	0x07, 0x32, 0x2D, 0x23, 0x50, 0x37, 0x3C, 0x08, 0x19, 0x59, 0x1F, 0x06,
	0x04, 0x47, 0x07, 0x08, 0x25, 0x15, 0x39, 0x0E, 0x1F, 0x03, 0x74, 0x02,
	0x03, 0x5B, 0x0C, 0x2C, 0x0F, 0x28, 0x5A, 0x5E, 0x29, 0x14, 0x57, 0x5C,
	0x29, 0x30, 0x38, 0x57, 0x36, 0x1B, 0x2C, 0x04, 0x28, 0x57, 0x09, 0x70,
	0x0E, 0x20, 0x58, 0x19, 0x0C, 0x5E, 0x30, 0x17, 0x2C, 0x2A, 0x16, 0x17,
	0x39, 0x2D, 0x29, 0x18, 0x2A, 0x00, 0x08, 0x76, 0x23, 0x4A, 0x16, 0x21,
	0x03, 0x59, 0x36, 0x04, 0x53, 0x26, 0x1C, 0x33, 0x2C, 0x32, 0x71, 0x01,
	0x17, 0x5F, 0x21, 0x15, 0x19, 0x00, 0x5F, 0x29, 0x37, 0x3F, 0x2A, 0x37,
	0x1B, 0x0A, 0x03, 0x26, 0x3E, 0x2F, 0x18, 0x1E, 0x19, 0x3F, 0x59, 0x29,
	0x0B, 0x0D, 0x03, 0x07, 0x23, 0x16, 0x4A, 0x3B, 0x07, 0x11, 0x00, 0x56,
	0x23, 0x22, 0x0A, 0x03, 0x17, 0x20, 0x1A, 0x08, 0x5D, 0x12, 0x03, 0x25,
	0x17, 0x35, 0x26, 0x23, 0x12, 0x2F, 0x27, 0x1B, 0x01, 0x1B, 0x13, 0x3A,
	0x26, 0x41, 0x19, 0x23, 0x25, 0x16, 0x5F, 0x20, 0x0C, 0x26, 0x0E, 0x5C,
	0x3D, 0x3A, 0x5D, 0x39, 0x03, 0x5A, 0x6D, 0x2E, 0x0E, 0x1E, 0x2F, 0x06,
	0x07, 0x30, 0x1A, 0x21, 0x23, 0x3A, 0x35, 0x01, 0x1A, 0x18, 0x23, 0x20,
	0x0B, 0x0E, 0x08, 0x5F, 0x51, 0x16, 0x1E, 0x23, 0x24, 0x50, 0x3E, 0x33,
	0x74, 0x3B, 0x53, 0x3A, 0x1A, 0x2E, 0x22, 0x00, 0x16, 0x28, 0x16, 0x15,
	0x10, 0x08, 0x3B, 0x2F, 0x22, 0x13, 0x27, 0x07, 0x2D, 0x1F, 0x53, 0x45,
	0x1B, 0x21, 0x39, 0x36, 0x5C, 0x39, 0x34, 0x5D, 0x0B, 0x0A, 0x09, 0x72,
	0x2B, 0x53, 0x39, 0x24, 0x38, 0x00, 0x55, 0x20, 0x5B, 0x25, 0x23, 0x53,
	0x3A, 0x3B, 0x33, 0x29, 0x52, 0x1A, 0x28, 0x13, 0x08, 0x00, 0x00, 0x32,
	0x23, 0x18, 0x27, 0x2C, 0x1D, 0x7B, 0x3D, 0x51, 0x1B, 0x1B, 0x09, 0x38,
	0x2A, 0x29, 0x05, 0x2D, 0x1D, 0x52, 0x00, 0x3B, 0x0C, 0x38, 0x58, 0x36,
	0x2F, 0x7B, 0x08, 0x57, 0x29, 0x52, 0x14, 0x27, 0x32, 0x0A, 0x44, 0x0E,
	0x22, 0x33, 0x39, 0x12, 0x08, 0x03, 0x13, 0x38, 0x5A, 0x75, 0x0A, 0x25,
	0x5F, 0x19, 0x00, 0x1A, 0x20, 0x3F, 0x5D, 0x74, 0x01, 0x0D, 0x07, 0x1B,
	0x08, 0x22, 0x17, 0x02, 0x07, 0x0B, 0x19, 0x07, 0x0F, 0x1D, 0x2D, 0x5C,
	0x17, 0x1C, 0x3A, 0x33, 0x59, 0x28, 0x05, 0x0F, 0x26, 0x2B, 0x57, 0x5B,
	0x13, 0x26, 0x36, 0x58, 0x1C, 0x44, 0x74, 0x22, 0x19, 0x0A, 0x1D, 0x73,
	0x26, 0x26, 0x3D, 0x02, 0x74, 0x25, 0x3B, 0x25, 0x1F, 0x20, 0x27, 0x00,
	0x5B, 0x1D, 0x10, 0x24, 0x10, 0x2D, 0x3A, 0x24, 0x0B, 0x33, 0x56, 0x05,
	0x76, 0x05, 0x33, 0x3A, 0x25, 0x13, 0x2A, 0x11, 0x06, 0x0A, 0x35, 0x3B,
	0x20, 0x1D, 0x1C, 0x31, 0x1E, 0x2D, 0x39, 0x5E, 0x71, 0x07, 0x29, 0x23,
	0x0C, 0x77, 0x5F, 0x35, 0x56, 0x12, 0x2D, 0x1D, 0x34, 0x57, 0x12, 0x37,
	0x3E, 0x56, 0x05, 0x03, 0x2B, 0x3F, 0x0B, 0x1A, 0x39, 0x11, 0x0E, 0x53,
	0x02, 0x3A, 0x18, 0x2E, 0x18, 0x5F, 0x33, 0x3B, 0x1A, 0x0C, 0x04, 0x59,
	0x32, 0x43, 0x4A, 0x22, 0x1B, 0x16, 0x09, 0x0E, 0x3D, 0x33, 0x29, 0x1B,
	0x53, 0x14, 0x0D, 0x29, 0x3E, 0x2E, 0x58, 0x3F, 0x0D, 0x55, 0x00, 0x00,
	0x01, 0x14, 0x01, 0x50, 0x1E, 0x5B, 0x7B, 0x2E, 0x57, 0x2A, 0x01, 0x37,
	0x18, 0x07, 0x1E, 0x1E, 0x73, 0x0F, 0x15, 0x21, 0x09, 0x06, 0x2A, 0x56,
	0x1B, 0x24, 0x25, 0x04, 0x10, 0x5F, 0x3E, 0x23, 0x18, 0x59, 0x27, 0x22,
	0x23, 0x1A, 0x00, 0x25, 0x0A, 0x36, 0x0D, 0x12, 0x23, 0x0F, 0x12, 0x09,
	0x39, 0x1A, 0x18, 0x1B, 0x27, 0x0F, 0x1E, 0x1A, 0x21, 0x18, 0x2A, 0x28,
	0x09, 0x18, 0x3E, 0x00, 0x16, 0x58, 0x2B, 0x0F, 0x35, 0x57, 0x1C, 0x2A,
	0x5E, 0x59, 0x06, 0x08, 0x16, 0x59, 0x07, 0x0A, 0x12, 0x76, 0x06, 0x15,
	0x2A, 0x52, 0x30, 0x35, 0x2E, 0x41, 0x1F, 0x27, 0x0D, 0x32, 0x06, 0x32,
	0x70, 0x5A, 0x19, 0x03, 0x26, 0x76, 0x04, 0x2F, 0x37, 0x5A, 0x26, 0x1E,
	0x28, 0x22, 0x5B, 0x21, 0x27, 0x14, 0x22, 0x25, 0x04, 0x26, 0x19, 0x04,
	0x38, 0x24, 0x0A, 0x06, 0x21, 0x01, 0x2C, 0x5A, 0x50, 0x23, 0x00, 0x0F,
	0x2A, 0x17, 0x36, 0x2D, 0x2B, 0x3F, 0x13, 0x1A, 0x03, 0x35, 0x18, 0x34,
	0x5E, 0x2E, 0x15, 0x29, 0x29, 0x27, 0x5A, 0x2B, 0x36, 0x4E, 0x5C, 0x3F,
	0x04, 0x3A, 0x02, 0x19, 0x07, 0x75, 0x3A, 0x00, 0x1A, 0x25, 0x25, 0x05,
	0x04, 0x5D, 0x3E, 0x35, 0x38, 0x31, 0x3D, 0x1F, 0x0F, 0x02, 0x53, 0x23,
	0x19, 0x77, 0x3B, 0x0E, 0x19, 0x1B, 0x77, 0x2B, 0x1B, 0x5B, 0x09, 0x14,
	0x16, 0x03, 0x2C, 0x2E, 0x7B, 0x00, 0x37, 0x1E, 0x24, 0x1B, 0x54, 0x31,
	0x1E, 0x39, 0x7B, 0x38, 0x19, 0x17, 0x2E, 0x18, 0x1E, 0x08, 0x5F, 0x38,
	0x0D, 0x3C, 0x30, 0x20, 0x03, 0x73, 0x3D, 0x0C, 0x08, 0x21, 0x72, 0x38,
	0x19, 0x57, 0x1A, 0x7B, 0x1A, 0x38, 0x5C, 0x3C, 0x2B, 0x07, 0x59, 0x34,
	0x44, 0x26, 0x1F, 0x17, 0x5B, 0x0C, 0x34, 0x00, 0x04, 0x18, 0x2E, 0x30,
	0x39, 0x2F, 0x5A, 0x0C, 0x16, 0x23, 0x15, 0x1B, 0x21, 0x33, 0x0F, 0x50,
	0x45, 0x25, 0x25, 0x14, 0x50, 0x5D, 0x5E, 0x08, 0x03, 0x29, 0x0F, 0x5E,
	0x2F, 0x3E, 0x0A, 0x56, 0x5F, 0x71, 0x3B, 0x37, 0x38, 0x21, 0x38, 0x2F,
	0x15, 0x0C, 0x27, 0x2B, 0x3A, 0x11, 0x45, 0x09, 0x0A, 0x2E, 0x17, 0x3C,
	0x40, 0x04, 0x21, 0x11, 0x5D, 0x32, 0x75, 0x24, 0x1B, 0x07, 0x25, 0x15,
	0x34, 0x37, 0x26, 0x25, 0x69, 0x06, 0x11, 0x3D, 0x19, 0x13, 0x5D, 0x0E,
	0x02, 0x01, 0x0C, 0x09, 0x06, 0x5D, 0x2E, 0x05, 0x55, 0x38, 0x0F, 0x3D,
	0x10, 0x1E, 0x50, 0x0D, 0x5F, 0x13, 0x59, 0x00, 0x1A, 0x2D, 0x04, 0x1A,
	0x0A, 0x57, 0x05, 0x0C, 0x19, 0x55, 0x38, 0x3E, 0x1A, 0x1E, 0x05, 0x3F,
	0x38, 0x70, 0x0D, 0x51, 0x5E, 0x32, 0x27, 0x0B, 0x04, 0x5F, 0x3F, 0x24,
	0x07, 0x32, 0x0D, 0x59, 0x2C, 0x34, 0x50, 0x04, 0x58, 0x76, 0x05, 0x2A,
	0x1F, 0x24, 0x33, 0x09, 0x53, 0x3D, 0x28, 0x14, 0x39, 0x25, 0x0D, 0x09,
	0x70, 0x00, 0x0C, 0x3C, 0x13, 0x2D, 0x5D, 0x4A, 0x56, 0x1F, 0x23, 0x1C,
	0x0A, 0x5C, 0x19, 0x32, 0x3A, 0x05, 0x01, 0x40, 0x28, 0x3E, 0x13, 0x1D,
	0x0A, 0x2F, 0x0A, 0x2E, 0x26, 0x3B, 0x1A, 0x15, 0x1B, 0x29, 0x38, 0x11,
	0x1D, 0x54, 0x0D, 0x33, 0x33, 0x00, 0x08, 0x1C, 0x5D, 0x11, 0x00, 0x2B,
	0x20, 0x22, 0x38, 0x02, 0x07, 0x0C, 0x18, 0x2A, 0x38, 0x2C, 0x5D, 0x05,
	0x27, 0x0B, 0x2E, 0x20, 0x1F, 0x13, 0x1A, 0x37, 0x16, 0x5A, 0x11, 0x3E,
	0x27, 0x2D, 0x0E, 0x28, 0x16, 0x20, 0x5E, 0x1D, 0x04, 0x54, 0x14, 0x2A,
	0x25, 0x0F, 0x5C, 0x55, 0x5A, 0x0E, 0x17, 0x5C, 0x02, 0x23, 0x19, 0x26,
	0x54, 0x24, 0x01, 0x5A, 0x72, 0x22, 0x39, 0x45, 0x32, 0x2B, 0x08, 0x10,
	0x1F, 0x52, 0x0C, 0x1C, 0x11, 0x2D, 0x44, 0x16, 0x36, 0x17, 0x5F, 0x03,
	0x7A, 0x55, 0x57, 0x0A, 0x19, 0x7B, 0x3E, 0x31, 0x3E, 0x24, 0x30, 0x55,
	0x00, 0x5F, 0x0E, 0x09, 0x14, 0x53, 0x3B, 0x19, 0x0E, 0x20, 0x05, 0x22,
	0x5F, 0x37, 0x19, 0x32, 0x23, 0x0A, 0x32, 0x0F, 0x33, 0x5D, 0x59, 0x6D,
	0x5B, 0x33, 0x1F, 0x25, 0x25, 0x00, 0x09, 0x5B, 0x07, 0x70, 0x35, 0x29,
	0x39, 0x0A, 0x0C, 0x5F, 0x20, 0x5D, 0x5A, 0x15, 0x19, 0x55, 0x2B, 0x59,
	0x01, 0x0A, 0x2E, 0x03, 0x5A, 0x2D, 0x2A, 0x37, 0x3A, 0x25, 0x11, 0x26,
	0x37, 0x34, 0x38, 0x2F, 0x5E, 0x0D, 0x16, 0x32, 0x76, 0x5A, 0x0A, 0x1D,
	0x11, 0x0F, 0x06, 0x04, 0x38, 0x5F, 0x2A, 0x3F, 0x17, 0x45, 0x32, 0x20,
	0x26, 0x16, 0x03, 0x12, 0x3B, 0x35, 0x57, 0x34, 0x2F, 0x30, 0x00, 0x2C,
	0x17, 0x1D, 0x2A, 0x23, 0x05, 0x57, 0x59, 0x18, 0x3F, 0x27, 0x27, 0x5A,
	0x06, 0x2E, 0x51, 0x20, 0x0A, 0x14, 0x0A, 0x0D, 0x1B, 0x3F, 0x27, 0x2A,
	0x0C, 0x5A, 0x20, 0x35, 0x2B, 0x37, 0x39, 0x1A, 0x12, 0x2E, 0x15, 0x2A,
	0x1F, 0x07, 0x55, 0x27, 0x0C, 0x33, 0x00, 0x2E, 0x13, 0x57, 0x5D, 0x70,
	0x21, 0x34, 0x05, 0x5A, 0x30, 0x1A, 0x39, 0x0B, 0x11, 0x72, 0x36, 0x3B,
	0x06, 0x5E, 0x0D, 0x3F, 0x36, 0x0F, 0x1F, 0x09, 0x28, 0x0D, 0x05, 0x52,
	0x05, 0x03, 0x09, 0x2A, 0x0E, 0x25, 0x1E, 0x04, 0x29, 0x07, 0x06, 0x07,
	0x00, 0x28, 0x18, 0x38, 0x1C, 0x31, 0x28, 0x2D, 0x0A, 0x16, 0x0B, 0x0A,
	0x5F, 0x7A, 0x2D, 0x03, 0x21, 0x3B, 0x35, 0x54, 0x03, 0x21, 0x58, 0x13,
	0x1D, 0x55, 0x19, 0x5B, 0x34, 0x0D, 0x58, 0x27, 0x3C, 0x36, 0x03, 0x51,
	0x0D, 0x0F, 0x34, 0x55, 0x00, 0x1F, 0x00, 0x23, 0x08, 0x2C, 0x21, 0x32,
	0x74, 0x3D, 0x32, 0x06, 0x2F, 0x36, 0x36, 0x30, 0x25, 0x59, 0x07, 0x15,
	0x37, 0x02, 0x40, 0x36, 0x1C, 0x18, 0x5F, 0x13, 0x00, 0x04, 0x0D, 0x5B,
	0x12, 0x23, 0x14, 0x25, 0x3F, 0x3A, 0x74, 0x55, 0x55, 0x25, 0x22, 0x06,
	0x0E, 0x35, 0x3A, 0x07, 0x3B, 0x24, 0x50, 0x27, 0x12, 0x2A, 0x47, 0x3B,
	0x1C, 0x13, 0x3A, 0x0F, 0x2B, 0x59, 0x13, 0x2E, 0x18, 0x1B, 0x5E, 0x31,
	0x75, 0x38, 0x2B, 0x01, 0x2E, 0x25, 0x15, 0x12, 0x5C, 0x1D, 0x13, 0x21,
	0x1B, 0x0A, 0x00, 0x38, 0x23, 0x53, 0x3F, 0x3E, 0x0D, 0x08, 0x57, 0x1F,
	0x12, 0x13, 0x2A, 0x2F, 0x2A, 0x28, 0x37, 0x38, 0x27, 0x0F, 0x2F, 0x2C,
	0x06, 0x26, 0x38, 0x21, 0x0A, 0x28, 0x3B, 0x20, 0x24, 0x2C, 0x26, 0x0B,
	0x23, 0x03, 0x28, 0x06, 0x2C, 0x5D, 0x24, 0x0C, 0x21, 0x50, 0x3A, 0x04,
	0x76, 0x08, 0x33, 0x3F, 0x12, 0x21, 0x03, 0x12, 0x23, 0x5E, 0x34, 0x16,
	0x0D, 0x2F, 0x5C, 0x15, 0x09, 0x18, 0x05, 0x5E, 0x03, 0x23, 0x0D, 0x5B,
	0x5D, 0x16, 0x34, 0x53, 0x57, 0x09, 0x35, 0x1B, 0x2C, 0x0B, 0x53, 0x2B,
	0x3A, 0x34, 0x3D, 0x26, 0x7A, 0x59, 0x2A, 0x04, 0x1F, 0x3A, 0x27, 0x0C,
	0x5D, 0x5B, 0x0C, 0x35, 0x56, 0x58, 0x44, 0x3B, 0x0A, 0x0A, 0x2D, 0x12,
	0x08, 0x22, 0x36, 0x03, 0x2F, 0x12, 0x21, 0x12, 0x16, 0x1D, 0x0A, 0x1A,
	0x15, 0x2D, 0x31, 0x37, 0x34, 0x08, 0x22, 0x0D, 0x2E, 0x22, 0x52, 0x56,
	0x13, 0x73, 0x02, 0x0D, 0x1E, 0x05, 0x04, 0x22, 0x13, 0x3B, 0x28, 0x3B,
	0x19, 0x57, 0x04, 0x33, 0x72, 0x20, 0x30, 0x3D, 0x0C, 0x33, 0x2B, 0x20,
	0x1B, 0x0D, 0x1B, 0x08, 0x0E, 0x1D, 0x5B, 0x74, 0x2B, 0x2A, 0x19, 0x33,
	0x29, 0x3A, 0x14, 0x0D, 0x03, 0x04, 0x1E, 0x37, 0x41, 0x3E, 0x35, 0x18,
	0x28, 0x29, 0x04, 0x75, 0x3D, 0x38, 0x38, 0x1B, 0x7B, 0x29, 0x00, 0x1D,
	0x21, 0x28, 0x5F, 0x08, 0x17, 0x2A, 0x74, 0x27, 0x0F, 0x03, 0x39, 0x74,
	0x1D, 0x09, 0x28, 0x52, 0x2E, 0x2B, 0x14, 0x25, 0x5A, 0x1A, 0x0D, 0x38,
	0x1D, 0x3F, 0x01, 0x1C, 0x20, 0x45, 0x09, 0x32, 0x24, 0x26, 0x21, 0x05,
	0x3A, 0x39, 0x2B, 0x3E, 0x59, 0x09, 0x27, 0x4A, 0x03, 0x18, 0x76, 0x27,
	0x29, 0x0A, 0x22, 0x00, 0x07, 0x4E, 0x18, 0x02, 0x35, 0x25, 0x07, 0x45,
	0x1E, 0x20, 0x43, 0x37, 0x29, 0x2D, 0x08, 0x19, 0x36, 0x14, 0x27, 0x0B,
	0x23, 0x34, 0x3A, 0x29, 0x34, 0x5A, 0x1B, 0x3D, 0x3C, 0x77, 0x5F, 0x12,
	0x14, 0x06, 0x00, 0x47, 0x34, 0x1C, 0x3B, 0x0F, 0x0D, 0x2D, 0x5F, 0x3C,
	0x0A, 0x1E, 0x16, 0x04, 0x19, 0x37, 0x54, 0x00, 0x0F, 0x5D, 0x21, 0x5C,
	0x0E, 0x2A, 0x04, 0x08, 0x09, 0x15, 0x1D, 0x5B, 0x77, 0x25, 0x53, 0x14,
	0x19, 0x16, 0x25, 0x07, 0x1A, 0x38, 0x05, 0x02, 0x2E, 0x5A, 0x3F, 0x15,
	0x23, 0x12, 0x1F, 0x40, 0x20, 0x20, 0x02, 0x1F, 0x05, 0x17, 0x21, 0x12,
	0x5D, 0x03, 0x34, 0x2E, 0x03, 0x22, 0x3A, 0x72, 0x0D, 0x24, 0x5D, 0x06,
	0x17, 0x36, 0x59, 0x0B, 0x1C, 0x2F, 0x36, 0x4E, 0x25, 0x06, 0x7B, 0x35,
	0x2B, 0x2B, 0x44, 0x09, 0x5E, 0x22, 0x1E, 0x04, 0x6D, 0x54, 0x37, 0x2A,
	0x2F, 0x20, 0x03, 0x50, 0x0D, 0x44, 0x2D, 0x3B, 0x14, 0x5D, 0x1A, 0x04,
	0x1A, 0x0C, 0x1F, 0x01, 0x05, 0x2F, 0x02, 0x1B, 0x27, 0x7A, 0x43, 0x04,
	0x17, 0x0E, 0x23, 0x1C, 0x38, 0x2F, 0x1F, 0x0C, 0x35, 0x28, 0x29, 0x11,
	0x36, 0x01, 0x22, 0x37, 0x11, 0x38, 0x22, 0x23, 0x09, 0x3B, 0x0C, 0x2A,
	0x10, 0x3B, 0x3D, 0x34, 0x2A, 0x29, 0x00, 0x40, 0x73, 0x26, 0x39, 0x5E,
	0x2E, 0x11, 0x03, 0x2D, 0x17, 0x20, 0x30, 0x1E, 0x00, 0x0F, 0x12, 0x32,
	0x00, 0x2C, 0x21, 0x2D, 0x34, 0x29, 0x22, 0x36, 0x32, 0x15, 0x5F, 0x1B,
	0x01, 0x02, 0x05, 0x1C, 0x00, 0x14, 0x5A, 0x2E, 0x5C, 0x08, 0x57, 0x52,
	0x2E, 0x0A, 0x56, 0x2F, 0x20, 0x29, 0x21, 0x13, 0x21, 0x07, 0x11, 0x07,
	0x13, 0x1D, 0x00, 0x15, 0x00, 0x28, 0x1E, 0x0A, 0x0C, 0x2A, 0x31, 0x14,
	0x3B, 0x09, 0x28, 0x11, 0x5C, 0x1B, 0x2A, 0x00, 0x13, 0x1E, 0x22, 0x16,
	0x21, 0x37, 0x24, 0x32, 0x25, 0x06, 0x23, 0x14, 0x1D, 0x0C, 0x20, 0x05,
	0x57, 0x26, 0x00, 0x3B, 0x12, 0x5C, 0x3F, 0x07, 0x15, 0x30, 0x1C, 0x0A,
	0x2D, 0x5D, 0x54, 0x25, 0x44, 0x38, 0x55, 0x56, 0x38, 0x02, 0x25, 0x5E,
	0x34, 0x37, 0x12, 0x1B, 0x18, 0x00, 0x2A, 0x3F, 0x23, 0x09, 0x1B, 0x5C,
	0x29, 0x6D, 0x21, 0x2E, 0x1C, 0x0A, 0x2E, 0x2E, 0x19, 0x07, 0x2D, 0x75,
	0x25, 0x24, 0x01, 0x2D, 0x72, 0x38, 0x12, 0x24, 0x12, 0x72, 0x02, 0x00,
	0x2B, 0x12, 0x6D, 0x36, 0x50, 0x0A, 0x06, 0x2E, 0x5B, 0x33, 0x04, 0x5C,
	0x26, 0x24, 0x28, 0x41, 0x0F, 0x1A, 0x15, 0x27, 0x1E, 0x59, 0x7B, 0x02,
	0x07, 0x04, 0x3A, 0x15, 0x3A, 0x10, 0x3B, 0x31, 0x08, 0x01, 0x4E, 0x27,
	0x29, 0x0C, 0x26, 0x35, 0x0A, 0x5A, 0x34, 0x5D, 0x15, 0x2D, 0x38, 0x03,
	0x03, 0x37, 0x38, 0x3B, 0x20, 0x5C, 0x09, 0x03, 0x0D, 0x20, 0x18, 0x00,
	0x1C, 0x38, 0x16, 0x22, 0x17, 0x22, 0x1C, 0x00, 0x01, 0x18, 0x41, 0x00,
	0x09, 0x1E, 0x15, 0x07, 0x3D, 0x09, 0x1C, 0x34, 0x14, 0x2C, 0x74, 0x35,
	0x33, 0x2D, 0x59, 0x2C, 0x25, 0x00, 0x22, 0x11, 0x26, 0x22, 0x12, 0x5A,
	0x01, 0x21, 0x3E, 0x3B, 0x39, 0x25, 0x24, 0x5E, 0x07, 0x28, 0x0A, 0x08,
	0x20, 0x06, 0x19, 0x25, 0x73, 0x07, 0x0A, 0x3A, 0x25, 0x0B, 0x36, 0x24,
	0x0D, 0x27, 0x06, 0x16, 0x32, 0x1E, 0x0A, 0x0F, 0x59, 0x05, 0x01, 0x1F,
	0x25, 0x14, 0x19, 0x0A, 0x38, 0x11, 0x26, 0x2E, 0x18, 0x24, 0x38, 0x05,
	0x2E, 0x1C, 0x5C, 0x01, 0x22, 0x05, 0x2D, 0x0F, 0x2F, 0x16, 0x0E, 0x3C,
	0x40, 0x75, 0x5D, 0x2D, 0x1D, 0x00, 0x37, 0x38, 0x2B, 0x28, 0x5D, 0x11,
	0x3C, 0x0D, 0x19, 0x3D, 0x1B, 0x5F, 0x32, 0x0C, 0x5A, 0x10, 0x5B, 0x32,
	0x24, 0x2A, 0x18, 0x18, 0x17, 0x5F, 0x21, 0x24, 0x19, 0x34, 0x23, 0x3C,
	0x2B, 0x36, 0x10, 0x18, 0x0F, 0x0F, 0x1C, 0x28, 0x01, 0x5D, 0x2E, 0x22,
	0x56, 0x29, 0x3A, 0x0E, 0x36, 0x51, 0x08, 0x25, 0x35, 0x03, 0x58, 0x29,
	0x28, 0x31, 0x47, 0x14, 0x57, 0x3C, 0x13, 0x29, 0x26, 0x05, 0x08, 0x24,
	0x5D, 0x04, 0x1C, 0x06, 0x72, 0x06, 0x50, 0x18, 0x0A, 0x36, 0x2F, 0x2C,
	0x1A, 0x2E, 0x34, 0x25, 0x2F, 0x19, 0x44, 0x17, 0x27, 0x56, 0x23, 0x59,
	0x25, 0x1E, 0x2C, 0x2F, 0x26, 0x38, 0x55, 0x33, 0x1C, 0x3C, 0x33, 0x07,
	0x15, 0x5F, 0x18, 0x2F, 0x1B, 0x26, 0x1A, 0x38, 0x14, 0x0A, 0x37, 0x58,
	0x04, 0x08, 0x18, 0x06, 0x16, 0x5C, 0x3B, 0x14, 0x2A, 0x03, 0x21, 0x04,
	0x03, 0x15, 0x14, 0x1F, 0x11, 0x28, 0x07, 0x2B, 0x1C, 0x74, 0x5B, 0x37,
	0x39, 0x12, 0x3B, 0x34, 0x29, 0x36, 0x52, 0x35, 0x1F, 0x37, 0x1C, 0x59,
	0x7A, 0x3E, 0x28, 0x1A, 0x3E, 0x33, 0x21, 0x10, 0x2A, 0x0E, 0x35, 0x00,
	0x11, 0x3B, 0x21, 0x05, 0x3B, 0x27, 0x16, 0x24, 0x29, 0x55, 0x56, 0x3A,
	0x12, 0x76, 0x3F, 0x2F, 0x3E, 0x05, 0x06, 0x07, 0x0A, 0x56, 0x21, 0x71,
	0x1E, 0x27, 0x1E, 0x32, 0x10, 0x47, 0x09, 0x17, 0x2C, 0x17, 0x58, 0x08,
	0x3D, 0x04, 0x24, 0x2F, 0x38, 0x1B, 0x0E, 0x38, 0x04, 0x51, 0x03, 0x31,
	0x2F, 0x38, 0x0E, 0x04, 0x05, 0x71, 0x5C, 0x22, 0x01, 0x5C, 0x72, 0x5A,
	0x04, 0x37, 0x2C, 0x0D, 0x3C, 0x32, 0x34, 0x26, 0x69, 0x54, 0x19, 0x57,
	0x24, 0x08, 0x5F, 0x53, 0x5B, 0x21, 0x2D, 0x1C, 0x15, 0x1F, 0x1C, 0x2B,
	0x35, 0x11, 0x58, 0x21, 0x18, 0x5D, 0x56, 0x57, 0x0A, 0x34, 0x26, 0x06,
	0x57, 0x0F, 0x38, 0x36, 0x2D, 0x22, 0x32, 0x28, 0x26, 0x4E, 0x1E, 0x0E,
	0x30, 0x1C, 0x33, 0x5A, 0x5E, 0x71, 0x28, 0x38, 0x16, 0x53, 0x17, 0x2F,
	0x35, 0x2F, 0x29, 0x07, 0x3B, 0x39, 0x59, 0x21, 0x20, 0x1A, 0x50, 0x05,
	0x22, 0x26, 0x3C, 0x55, 0x0C, 0x3D, 0x27, 0x1C, 0x05, 0x23, 0x02, 0x04,
	0x27, 0x50, 0x21, 0x05, 0x11, 0x3F, 0x04, 0x1A, 0x31, 0x23, 0x3D, 0x3B,
	0x02, 0x32, 0x0B, 0x5A, 0x04, 0x17, 0x3B, 0x0D, 0x5D, 0x19, 0x45, 0x1E,
	0x73, 0x0F, 0x11, 0x02, 0x27, 0x73, 0x27, 0x17, 0x09, 0x1B, 0x31, 0x5C,
	0x20, 0x34, 0x1A, 0x13, 0x5D, 0x51, 0x1E, 0x0F, 0x0E, 0x0D, 0x29, 0x2A,
	0x2A, 0x2D, 0x2B, 0x58, 0x18, 0x5F, 0x74, 0x3E, 0x22, 0x06, 0x25, 0x2F,
	0x08, 0x27, 0x56, 0x2F, 0x16, 0x0A, 0x58, 0x05, 0x22, 0x0C, 0x3A, 0x3B,
	0x2A, 0x5F, 0x73, 0x3B, 0x3B, 0x0D, 0x06, 0x7A, 0x3F, 0x13, 0x18, 0x5B,
	0x35, 0x58, 0x12, 0x17, 0x09, 0x12, 0x07, 0x39, 0x38, 0x23, 0x09, 0x29,
	0x2C, 0x3D, 0x11, 0x3A, 0x16, 0x0D, 0x01, 0x03, 0x38, 0x43, 0x2D, 0x28,
	0x02, 0x0B, 0x3B, 0x11, 0x3D, 0x09, 0x34, 0x0E, 0x54, 0x04, 0x40, 0x77,
	0x1D, 0x3B, 0x17, 0x06, 0x08, 0x58, 0x0B, 0x3D, 0x25, 0x38, 0x36, 0x2A,
	0x5F, 0x33, 0x13, 0x34, 0x2F, 0x28, 0x07, 0x09, 0x2A, 0x53, 0x5B, 0x27,
	0x36, 0x54, 0x57, 0x5E, 0x5D, 0x74, 0x1D, 0x06, 0x17, 0x04, 0x2B, 0x19,
	0x0A, 0x24, 0x18, 0x0E, 0x01, 0x3B, 0x07, 0x12, 0x09, 0x07, 0x39, 0x27,
	0x5C, 0x09, 0x5E, 0x32, 0x39, 0x3F, 0x09, 0x06, 0x56, 0x39, 0x39, 0x70,
	0x3A, 0x19, 0x19, 0x11, 0x23, 0x01, 0x50, 0x1E, 0x3C, 0x7B, 0x54, 0x2C,
	0x1B, 0x0D, 0x77, 0x27, 0x2E, 0x34, 0x59, 0x13, 0x5A, 0x34, 0x2B, 0x02,
	0x04, 0x35, 0x28, 0x01, 0x0F, 0x0E, 0x15, 0x51, 0x36, 0x1E, 0x25, 0x22,
	0x08, 0x5A, 0x26, 0x13, 0x1B, 0x2B, 0x39, 0x52, 0x26, 0x54, 0x56, 0x1D,
	0x31, 0x0B, 0x3B, 0x15, 0x39, 0x2D, 0x1B, 0x2A, 0x0E, 0x1B, 0x3A, 0x09,
	0x1F, 0x52, 0x58, 0x27, 0x3A, 0x04, 0x05, 0x18, 0x00, 0x3B, 0x54, 0x4A,
	0x03, 0x24, 0x10, 0x14, 0x14, 0x1A, 0x07, 0x0C, 0x06, 0x09, 0x1B, 0x38,
	0x2C, 0x0E, 0x0F, 0x3D, 0x0E, 0x1B, 0x47, 0x0A, 0x04, 0x1A, 0x69, 0x0D,
	0x12, 0x2C, 0x12, 0x16, 0x20, 0x57, 0x3F, 0x5E, 0x36, 0x00, 0x06, 0x5D,
	0x21, 0x1B, 0x58, 0x12, 0x39, 0x3C, 0x69, 0x06, 0x34, 0x3C, 0x3E, 0x2F,
	0x07, 0x2C, 0x1E, 0x12, 0x18, 0x2B, 0x39, 0x0F, 0x08, 0x10, 0x55, 0x58,
	0x5A, 0x04, 0x29, 0x02, 0x39, 0x3D, 0x23, 0x06, 0x23, 0x25, 0x24, 0x21,
	0x17, 0x38, 0x0E, 0x39, 0x2C, 0x28, 0x3B, 0x57, 0x5B, 0x53, 0x3A, 0x25,
	0x30, 0x01, 0x3D, 0x06, 0x0D, 0x17, 0x45, 0x24, 0x1A, 0x0F, 0x35, 0x07,
	0x03, 0x15, 0x5D, 0x36, 0x1E, 0x33, 0x70, 0x0F, 0x1B, 0x1D, 0x3B, 0x18,
	0x1E, 0x2A, 0x03, 0x52, 0x01, 0x26, 0x3B, 0x07, 0x1C, 0x08, 0x01, 0x34,
	0x1E, 0x28, 0x0F, 0x16, 0x56, 0x26, 0x5D, 0x27, 0x34, 0x51, 0x5F, 0x1E,
	0x13, 0x2E, 0x2A, 0x28, 0x5A, 0x05, 0x1C, 0x27, 0x22, 0x5E, 0x07, 0x00,
	0x56, 0x59, 0x2C, 0x0A, 0x22, 0x2D, 0x5B, 0x24, 0x0E, 0x24, 0x02, 0x03,
	0x32, 0x12, 0x0E, 0x25, 0x39, 0x5D, 0x32, 0x3F, 0x08, 0x2C, 0x06, 0x11,
	0x03, 0x54, 0x0F, 0x08, 0x75, 0x20, 0x35, 0x3A, 0x20, 0x2C, 0x2D, 0x1B,
	0x36, 0x11, 0x37, 0x39, 0x2A, 0x3B, 0x0C, 0x75, 0x25, 0x28, 0x0B, 0x24,
	0x14, 0x28, 0x0B, 0x1B, 0x44, 0x0E, 0x0F, 0x11, 0x39, 0x21, 0x26, 0x36,
	0x53, 0x14, 0x3F, 0x36, 0x27, 0x25, 0x2B, 0x11, 0x0D, 0x3D, 0x00, 0x04,
	0x04, 0x38, 0x36, 0x39, 0x38, 0x22, 0x34, 0x55, 0x0A, 0x08, 0x2D, 0x2A,
	0x21, 0x2A, 0x20, 0x3C, 0x69, 0x3D, 0x2F, 0x1B, 0x0A, 0x30, 0x28, 0x57,
	0x07, 0x20, 0x12, 0x3C, 0x50, 0x23, 0x31, 0x28, 0x08, 0x24, 0x0B, 0x0D,
	0x71, 0x3F, 0x07, 0x00, 0x11, 0x0C, 0x47, 0x57, 0x41, 0x00, 0x29, 0x00,
	0x36, 0x0F, 0x59, 0x16, 0x3B, 0x04, 0x2C, 0x1E, 0x77, 0x2B, 0x2A, 0x09,
	0x5B, 0x11, 0x0E, 0x0F, 0x0D, 0x00, 0x01, 0x1A, 0x07, 0x3B, 0x2D, 0x76,
	0x27, 0x16, 0x00, 0x5D, 0x2F, 0x0E, 0x51, 0x18, 0x0F, 0x0A, 0x43, 0x15,
	0x3B, 0x00, 0x38, 0x38, 0x04, 0x21, 0x22, 0x28, 0x5C, 0x38, 0x3A, 0x33,
	0x33, 0x5D, 0x19, 0x3B, 0x39, 0x26, 0x47, 0x14, 0x3C, 0x58, 0x30, 0x47,
	0x1B, 0x2B, 0x03, 0x25, 0x29, 0x09, 0x05, 0x13, 0x2F, 0x00, 0x16, 0x26,
	0x09, 0x2A, 0x1B, 0x15, 0x1E, 0x06, 0x12, 0x18, 0x00, 0x0A, 0x3E, 0x27,
	0x22, 0x0F, 0x24, 0x28, 0x12, 0x55, 0x1B, 0x2A, 0x1F, 0x3A, 0x14, 0x50,
	0x17, 0x29, 0x34, 0x00, 0x0F, 0x26, 0x2F, 0x00, 0x1B, 0x2C, 0x18, 0x26,
	0x29, 0x39, 0x52, 0x37, 0x26, 0x06, 0x29, 0x16, 0x14, 0x18, 0x33, 0x5E,
	0x12, 0x3C, 0x5C, 0x33, 0x1C, 0x14, 0x5C, 0x5F, 0x30, 0x5D, 0x17, 0x34,
	0x1F, 0x1A, 0x36, 0x3B, 0x3B, 0x2C, 0x10, 0x09, 0x18, 0x3E, 0x0C, 0x2D,
	0x1D, 0x36, 0x0C, 0x22, 0x28, 0x38, 0x2D, 0x3C, 0x3F, 0x2D, 0x58, 0x51,
	0x03, 0x04, 0x3A, 0x00, 0x28, 0x57, 0x2C, 0x2C, 0x0A, 0x36, 0x45, 0x24,
	0x0C, 0x05, 0x3B, 0x34, 0x18, 0x05, 0x01, 0x11, 0x29, 0x1E, 0x76, 0x43,
	0x32, 0x0A, 0x59, 0x2A, 0x06, 0x12, 0x36, 0x03, 0x26, 0x2D, 0x22, 0x07,
	0x11, 0x30, 0x23, 0x51, 0x36, 0x0E, 0x7B, 0x38, 0x4E, 0x17, 0x5A, 0x3A,
	0x02, 0x50, 0x27, 0x5C, 0x38, 0x24, 0x39, 0x17, 0x19, 0x38, 0x35, 0x57,
	0x1A, 0x27, 0x32, 0x22, 0x37, 0x56, 0x1B, 0x31, 0x54, 0x2F, 0x1A, 0x0A,
	0x11, 0x08, 0x13, 0x19, 0x3E, 0x2B, 0x07, 0x54, 0x1B, 0x02, 0x3B, 0x39,
	0x15, 0x1A, 0x1F, 0x76, 0x1E, 0x14, 0x00, 0x0C, 0x3A, 0x36, 0x12, 0x2B,
	0x0D, 0x2A, 0x34, 0x24, 0x3B, 0x13, 0x14, 0x1D, 0x05, 0x2B, 0x08, 0x7B,
	0x1E, 0x52, 0x5C, 0x1A, 0x23, 0x3F, 0x54, 0x5D, 0x5A, 0x25, 0x20, 0x4A,
	0x45, 0x31, 0x17, 0x0F, 0x2C, 0x26, 0x0A, 0x7A, 0x0F, 0x0F, 0x3D, 0x3E,
	0x0D, 0x0D, 0x4E, 0x5C, 0x09, 0x07, 0x35, 0x57, 0x07, 0x26, 0x76, 0x5F,
	0x13, 0x28, 0x09, 0x1B, 0x25, 0x0F, 0x39, 0x0A, 0x38, 0x2F, 0x22, 0x26,
	0x22, 0x3B, 0x26, 0x55, 0x5B, 0x3A, 0x15, 0x0D, 0x2D, 0x1A, 0x25, 0x33,
	0x0D, 0x12, 0x03, 0x02, 0x25, 0x5E, 0x17, 0x34, 0x31, 0x11, 0x47, 0x50,
	0x03, 0x2D, 0x26, 0x05, 0x24, 0x45, 0x2F, 0x32, 0x28, 0x59, 0x24, 0x2D,
	0x31, 0x26, 0x2E, 0x59, 0x3C, 0x25, 0x14, 0x2B, 0x5F, 0x5B, 0x28, 0x20,
	0x25, 0x36, 0x32, 0x70, 0x58, 0x55, 0x16, 0x40, 0x33, 0x21, 0x2A, 0x2B,
	0x0D, 0x0A, 0x1A, 0x3B, 0x39, 0x5D, 0x25, 0x16, 0x30, 0x03, 0x06, 0x04,
	0x14, 0x3B, 0x16, 0x3A, 0x06, 0x25, 0x14, 0x3B, 0x22, 0x77, 0x3A, 0x2C,
	0x0A, 0x04, 0x35, 0x00, 0x50, 0x37, 0x44, 0x16, 0x3A, 0x24, 0x2F, 0x05,
	0x37, 0x1C, 0x02, 0x0A, 0x20, 0x32, 0x03, 0x54, 0x24, 0x5A, 0x2E, 0x39,
	0x22, 0x5B, 0x3B, 0x69, 0x1C, 0x55, 0x5C, 0x24, 0x17, 0x2F, 0x50, 0x08,
	0x5D, 0x13, 0x1C, 0x10, 0x1B, 0x22, 0x07, 0x1A, 0x25, 0x39, 0x32, 0x2C,
	0x58, 0x51, 0x01, 0x1F, 0x06, 0x22, 0x08, 0x02, 0x03, 0x2C, 0x38, 0x03,
	0x1C, 0x24, 0x12, 0x3B, 0x15, 0x5A, 0x33, 0x01, 0x3A, 0x32, 0x39, 0x24,
	0x3A, 0x34, 0x55, 0x3E, 0x5C, 0x10, 0x35, 0x0A, 0x3F, 0x31, 0x38, 0x19,
	0x37, 0x2A, 0x01, 0x18, 0x28, 0x53, 0x08, 0x12, 0x01, 0x3F, 0x17, 0x0B,
	0x22, 0x32, 0x0F, 0x03, 0x5A, 0x3C, 0x1B, 0x3E, 0x03, 0x08, 0x0C, 0x2E,
	0x2A, 0x19, 0x56, 0x26, 0x29, 0x19, 0x51, 0x19, 0x1B, 0x2C, 0x47, 0x0C,
	0x58, 0x52, 0x1B, 0x01, 0x52, 0x23, 0x0F, 0x12, 0x1D, 0x29, 0x08, 0x23,
	0x0D, 0x3E, 0x0E, 0x58, 0x08, 0x18, 0x03, 0x1B, 0x0C, 0x2A, 0x2B, 0x3A,
	0x10, 0x45, 0x32, 0x2C, 0x28, 0x11, 0x1A, 0x2F, 0x2E, 0x2A, 0x37, 0x5F,
	0x24, 0x09, 0x1F, 0x32, 0x5C, 0x25, 0x0A, 0x1D, 0x0A, 0x22, 0x1A, 0x11,
	0x26, 0x2C, 0x3A, 0x31, 0x12, 0x34, 0x11, 0x05, 0x2A, 0x24, 0x3D, 0x13,
	0x3B, 0x5B, 0x0F, 0x2A, 0x36, 0x3B, 0x12, 0x27, 0x3B, 0x2D, 0x02, 0x0A,
	0x14, 0x0F, 0x27, 0x58, 0x5F, 0x2D, 0x5A, 0x0E, 0x22, 0x11, 0x2A, 0x38,
	0x25, 0x3C, 0x1E, 0x08, 0x24, 0x30, 0x3E, 0x58, 0x71, 0x26, 0x0D, 0x23,
	0x03, 0x0B, 0x04, 0x1B, 0x02, 0x0E, 0x70, 0x5C, 0x55, 0x3F, 0x39, 0x07,
	0x02, 0x31, 0x3B, 0x25, 0x71, 0x05, 0x0B, 0x00, 0x19, 0x05, 0x59, 0x06,
	0x3C, 0x2F, 0x31, 0x5B, 0x4A, 0x0D, 0x07, 0x18, 0x2F, 0x1B, 0x3A, 0x1D,
	0x17, 0x36, 0x33, 0x3F, 0x24, 0x27, 0x47, 0x08, 0x2A, 0x3B, 0x00, 0x47,
	0x58, 0x2D, 0x3F, 0x23, 0x25, 0x00, 0x3E, 0x2F, 0x26, 0x02, 0x25, 0x37,
	0x22, 0x69, 0x3C, 0x17, 0x59, 0x53, 0x35, 0x27, 0x0F, 0x3A, 0x3E, 0x20,
	0x38, 0x37, 0x20, 0x01, 0x3A, 0x38, 0x07, 0x59, 0x2C, 0x34, 0x3B, 0x0A,
	0x20, 0x21, 0x10, 0x0D, 0x11, 0x3D, 0x05, 0x05, 0x0E, 0x15, 0x58, 0x5B,
	0x69, 0x16, 0x06, 0x0A, 0x28, 0x37, 0x54, 0x0A, 0x19, 0x3C, 0x01, 0x18,
	0x2B, 0x2C, 0x1B, 0x31, 0x35, 0x00, 0x0D, 0x5D, 0x27, 0x5B, 0x29, 0x24,
	0x24, 0x2C, 0x2B, 0x32, 0x57, 0x0A, 0x29, 0x28, 0x18, 0x39, 0x5B, 0x09,
	0x1F, 0x37, 0x07, 0x0E, 0x38, 0x3A, 0x19, 0x08, 0x00, 0x1A, 0x18, 0x2D,
	0x0A, 0x26, 0x0B, 0x28, 0x2D, 0x5F, 0x24, 0x33, 0x19, 0x0D, 0x5A, 0x27,
	0x05, 0x54, 0x50, 0x06, 0x00, 0x77, 0x38, 0x10, 0x2C, 0x05, 0x09, 0x05,
	0x35, 0x0F, 0x5B, 0x76, 0x54, 0x3B, 0x0C, 0x06, 0x37, 0x5B, 0x2C, 0x17,
	0x21, 0x0C, 0x06, 0x3B, 0x2B, 0x22, 0x18, 0x0F, 0x25, 0x07, 0x06, 0x33,
	0x24, 0x10, 0x0F, 0x1A, 0x00, 0x27, 0x0B, 0x3B, 0x3A, 0x2B, 0x55, 0x57,
	0x28, 0x22, 0x2C, 0x04, 0x0D, 0x39, 0x09, 0x12, 0x54, 0x39, 0x1C, 0x08,
	0x04, 0x3A, 0x19, 0x56, 0x3F, 0x0C, 0x43, 0x35, 0x2B, 0x1A, 0x21, 0x07,
	0x39, 0x05, 0x01, 0x24, 0x20, 0x11, 0x05, 0x3E, 0x14, 0x0A, 0x05, 0x5C,
	0x53, 0x72, 0x43, 0x34, 0x0A, 0x3E, 0x25, 0x28, 0x26, 0x17, 0x40, 0x0B,
	0x1F, 0x54, 0x3C, 0x26, 0x12, 0x5A, 0x16, 0x20, 0x24, 0x69, 0x34, 0x14,
	0x25, 0x00, 0x77, 0x59, 0x59, 0x14, 0x2F, 0x16, 0x3F, 0x34, 0x16, 0x58,
	0x23, 0x3F, 0x36, 0x02, 0x0D, 0x36, 0x1B, 0x30, 0x0B, 0x21, 0x33, 0x1E,
	0x00, 0x06, 0x31, 0x03, 0x08, 0x33, 0x58, 0x08, 0x12, 0x5C, 0x29, 0x38,
	0x3A, 0x7A, 0x58, 0x33, 0x0F, 0x26, 0x2D, 0x09, 0x0F, 0x39, 0x2C, 0x07,
	0x01, 0x09, 0x3F, 0x23, 0x06, 0x19, 0x2B, 0x19, 0x5D, 0x2D, 0x2B, 0x1B,
	0x1D, 0x5B, 0x2E, 0x00, 0x04, 0x00, 0x21, 0x05, 0x5B, 0x54, 0x01, 0x39,
	0x71, 0x01, 0x16, 0x5D, 0x1F, 0x14, 0x0B, 0x53, 0x18, 0x53, 0x24, 0x35,
	0x33, 0x25, 0x25, 0x20, 0x04, 0x10, 0x5D, 0x3A, 0x01, 0x3E, 0x2E, 0x20,
	0x25, 0x2F, 0x0F, 0x0D, 0x58, 0x0D, 0x3A, 0x26, 0x2E, 0x1F, 0x3F, 0x69,
	0x55, 0x08, 0x27, 0x58, 0x26, 0x0D, 0x32, 0x28, 0x1D, 0x1B, 0x15, 0x51,
	0x0B, 0x1B, 0x73, 0x3C, 0x56, 0x29, 0x03, 0x0F, 0x34, 0x09, 0x14, 0x18,
	0x0F, 0x22, 0x34, 0x05, 0x32, 0x16, 0x2B, 0x37, 0x09, 0x5C, 0x2F, 0x0B,
	0x3B, 0x0D, 0x1A, 0x07, 0x3B, 0x25, 0x39, 0x01, 0x20, 0x39, 0x39, 0x1E,
	0x09, 0x73, 0x5D, 0x35, 0x0C, 0x2D, 0x14, 0x58, 0x39, 0x23, 0x52, 0x1A,
	0x34, 0x08, 0x5D, 0x1D, 0x0A, 0x09, 0x2B, 0x27, 0x28, 0x06, 0x01, 0x57,
	0x06, 0x0A, 0x01, 0x43, 0x3B, 0x1C, 0x1B, 0x1B, 0x5C, 0x0D, 0x36, 0x5F,
	0x31, 0x22, 0x15, 0x5E, 0x2D, 0x1A, 0x0B, 0x27, 0x18, 0x38, 0x20, 0x08,
	0x57, 0x3B, 0x0A, 0x34, 0x05, 0x35, 0x2A, 0x20, 0x15, 0x1C, 0x12, 0x59,
	0x1A, 0x10, 0x18, 0x37, 0x05, 0x28, 0x35, 0x2D, 0x2A, 0x24, 0x1D, 0x27,
	0x23, 0x27, 0x3D, 0x25, 0x18, 0x07, 0x29, 0x02, 0x58, 0x33, 0x1B, 0x2C,
	0x39, 0x59, 0x2D, 0x5A, 0x11, 0x57, 0x2D, 0x6D, 0x3E, 0x32, 0x18, 0x08,
	0x73, 0x2F, 0x3B, 0x5F, 0x3B, 0x08, 0x14, 0x51, 0x3F, 0x04, 0x75, 0x21,
	0x58, 0x27, 0x09, 0x3A, 0x39, 0x26, 0x04, 0x3C, 0x0C, 0x36, 0x2B, 0x5E,
	0x2D, 0x32, 0x34, 0x31, 0x29, 0x31, 0x23, 0x08, 0x33, 0x5D, 0x2A, 0x05,
	0x38, 0x15, 0x27, 0x39, 0x04, 0x58, 0x34, 0x02, 0x3E, 0x7B, 0x28, 0x39,
	0x36, 0x25, 0x03, 0x1F, 0x34, 0x22, 0x2F, 0x74, 0x26, 0x0D, 0x3E, 0x2E,
	0x28, 0x05, 0x05, 0x18, 0x09, 0x72, 0x2B, 0x26, 0x28, 0x06, 0x3B, 0x3D,
	0x19, 0x0A, 0x03, 0x1A, 0x59, 0x05, 0x07, 0x1A, 0x38, 0x0B, 0x0A, 0x34,
	0x04, 0x31, 0x54, 0x19, 0x3E, 0x0D, 0x00, 0x1D, 0x51, 0x25, 0x1E, 0x26,
	0x19, 0x05, 0x23, 0x23, 0x27, 0x2A, 0x0C, 0x38, 0x1B, 0x2D, 0x06, 0x4A,
	0x3B, 0x18, 0x2F, 0x08, 0x56, 0x01, 0x21, 0x33, 0x20, 0x2F, 0x20, 0x44,
	0x18, 0x1D, 0x39, 0x08, 0x3A, 0x2A, 0x5D, 0x14, 0x24, 0x20, 0x71, 0x3A,
	0x36, 0x0D, 0x05, 0x2D, 0x38, 0x53, 0x0D, 0x38, 0x3A, 0x5B, 0x05, 0x19,
	0x3D, 0x0B, 0x3C, 0x56, 0x16, 0x3F, 0x0B, 0x1F, 0x0B, 0x57, 0x2C, 0x0A,
	0x3E, 0x3B, 0x23, 0x08, 0x70, 0x1F, 0x22, 0x0D, 0x0F, 0x37, 0x28, 0x39,
	0x34, 0x23, 0x0C, 0x21, 0x20, 0x1F, 0x1E, 0x72, 0x43, 0x29, 0x2C, 0x33,
	0x15, 0x2F, 0x51, 0x5C, 0x04, 0x3B, 0x3F, 0x50, 0x3E, 0x08, 0x14, 0x22,
	0x2A, 0x03, 0x05, 0x05, 0x19, 0x0D, 0x17, 0x00, 0x2E, 0x25, 0x2C, 0x3A,
	0x38, 0x75, 0x2A, 0x07, 0x3C, 0x5D, 0x10, 0x3E, 0x08, 0x41, 0x12, 0x26,
	0x5E, 0x32, 0x1C, 0x58, 0x16, 0x1D, 0x36, 0x23, 0x1B, 0x05, 0x18, 0x0D,
	0x17, 0x1B, 0x72, 0x16, 0x34, 0x0D, 0x59, 0x14, 0x55, 0x23, 0x2C, 0x18,
	0x2D, 0x26, 0x33, 0x38, 0x19, 0x0C, 0x55, 0x54, 0x59, 0x5C, 0x38, 0x2D,
	0x03, 0x0B, 0x1A, 0x24, 0x01, 0x37, 0x3B, 0x08, 0x26, 0x0D, 0x35, 0x5F,
	0x00, 0x2E, 0x2A, 0x2A, 0x19, 0x02, 0x16, 0x36, 0x31, 0x1A, 0x04, 0x00,
	0x58, 0x35, 0x3F, 0x29, 0x0A, 0x3F, 0x10, 0x1A, 0x18, 0x27, 0x43, 0x2F,
	0x1C, 0x52, 0x73, 0x2B, 0x03, 0x14, 0x27, 0x7B, 0x07, 0x10, 0x3F, 0x2E,
	0x25, 0x02, 0x58, 0x56, 0x0C, 0x26, 0x1D, 0x59, 0x22, 0x31, 0x0D, 0x14,
	0x57, 0x5B, 0x3E, 0x29, 0x2E, 0x18, 0x07, 0x1B, 0x27, 0x54, 0x0F, 0x2C,
	0x21, 0x75, 0x34, 0x22, 0x5E, 0x13, 0x2D, 0x14, 0x30, 0x57, 0x25, 0x71,
	0x25, 0x09, 0x3E, 0x01, 0x0F, 0x18, 0x0F, 0x5B, 0x38, 0x72, 0x2F, 0x32,
	0x05, 0x13, 0x3A, 0x00, 0x03, 0x19, 0x1A, 0x03, 0x35, 0x51, 0x2B, 0x38,
	0x20, 0x5C, 0x38, 0x05, 0x07, 0x36, 0x05, 0x16, 0x34, 0x3C, 0x09, 0x36,
	0x08, 0x57, 0x03, 0x08, 0x1D, 0x57, 0x56, 0x5B, 0x27, 0x43, 0x03, 0x1D,
	0x12, 0x72, 0x3D, 0x0C, 0x1F, 0x59, 0x36, 0x02, 0x53, 0x02, 0x33, 0x2B,
	0x5E, 0x2E, 0x19, 0x00, 0x72, 0x34, 0x37, 0x19, 0x52, 0x1A, 0x0E, 0x39,
	0x20, 0x29, 0x17, 0x01, 0x1B, 0x3C, 0x39, 0x72, 0x1E, 0x25, 0x34, 0x52,
	0x0A, 0x5C, 0x3B, 0x21, 0x3F, 0x0F, 0x03, 0x08, 0x08, 0x20, 0x0B, 0x5E,
	0x2B, 0x5B, 0x00, 0x7B, 0x0B, 0x4A, 0x58, 0x26, 0x1B, 0x20, 0x28, 0x1F,
	0x39, 0x12, 0x21, 0x13, 0x5E, 0x1A, 0x17, 0x2B, 0x02, 0x5A, 0x38, 0x37,
	0x43, 0x06, 0x3B, 0x11, 0x71, 0x1F, 0x34, 0x1F, 0x32, 0x33, 0x18, 0x38,
	0x1F, 0x0A, 0x20, 0x38, 0x0B, 0x57, 0x2E, 0x2E, 0x3A, 0x12, 0x0B, 0x58,
	0x70, 0x03, 0x0F, 0x3E, 0x11, 0x03, 0x43, 0x2A, 0x0F, 0x5B, 0x07, 0x5E,
	0x2E, 0x0D, 0x03, 0x26, 0x5E, 0x03, 0x2D, 0x5C, 0x0B, 0x18, 0x52, 0x0D,
	0x39, 0x33, 0x1A, 0x15, 0x5C, 0x25, 0x1A, 0x19, 0x23, 0x1B, 0x1D, 0x0C,
	0x09, 0x33, 0x38, 0x18, 0x0F, 0x24, 0x2B, 0x24, 0x2C, 0x70, 0x47, 0x50,
	0x20, 0x19, 0x36, 0x39, 0x0B, 0x5F, 0x1C, 0x11, 0x2F, 0x2E, 0x16, 0x59,
	0x0C, 0x05, 0x4E, 0x2D, 0x27, 0x3A, 0x20, 0x1B, 0x1A, 0x20, 0x20, 0x07,
	0x2E, 0x29, 0x07, 0x11, 0x3A, 0x12, 0x28, 0x21, 0x70, 0x39, 0x19, 0x56,
	0x23, 0x04, 0x09, 0x15, 0x58, 0x33, 0x35, 0x38, 0x31, 0x45, 0x2C, 0x70,
	0x27, 0x50, 0x02, 0x38, 0x20, 0x47, 0x0C, 0x2B, 0x3D, 0x32, 0x5E, 0x14,
	0x34, 0x0F, 0x21, 0x2F, 0x58, 0x27, 0x31, 0x28, 0x2A, 0x04, 0x14, 0x06,
	0x20, 0x29, 0x50, 0x27, 0x21, 0x29, 0x07, 0x0C, 0x25, 0x19, 0x6D, 0x15,
	0x06, 0x28, 0x27, 0x70, 0x24, 0x07, 0x0C, 0x23, 0x6D, 0x0A, 0x4A, 0x1A,
	0x18, 0x32, 0x0D, 0x37, 0x24, 0x22, 0x2D, 0x26, 0x22, 0x1B, 0x0E, 0x73,
	0x39, 0x58, 0x06, 0x3E, 0x0E, 0x26, 0x33, 0x2C, 0x04, 0x71, 0x38, 0x2D,
	0x1C, 0x39, 0x72, 0x22, 0x15, 0x06, 0x22, 0x07, 0x16, 0x03, 0x2B, 0x1A,
	0x12, 0x38, 0x32, 0x24, 0x1D, 0x33, 0x38, 0x0B, 0x1E, 0x1F, 0x09, 0x08,
	0x26, 0x07, 0x29, 0x08, 0x58, 0x11, 0x3F, 0x24, 0x2D, 0x1F, 0x1B, 0x3E,
	0x58, 0x08, 0x39, 0x03, 0x0C, 0x11, 0x0A, 0x01, 0x14, 0x18, 0x1F, 0x08,
	0x3A, 0x22, 0x1F, 0x18, 0x28, 0x2A, 0x4A, 0x01, 0x27, 0x0B, 0x2E, 0x53,
	0x3A, 0x3E, 0x71, 0x26, 0x0A, 0x38, 0x06, 0x34, 0x5D, 0x12, 0x20, 0x2C,
	0x2F, 0x22, 0x06, 0x56, 0x11, 0x26, 0x1D, 0x36, 0x05, 0x08, 0x3A, 0x55,
	0x58, 0x3C, 0x26, 0x2B, 0x3E, 0x52, 0x5E, 0x0D, 0x28, 0x1C, 0x4E, 0x1A,
	0x09, 0x3A, 0x20, 0x13, 0x37, 0x2D, 0x70, 0x1E, 0x2F, 0x0A, 0x5B, 0x03,
	0x29, 0x0F, 0x03, 0x3D, 0x28, 0x18, 0x05, 0x57, 0x27, 0x15, 0x1E, 0x39,
	0x05, 0x01, 0x25, 0x1D, 0x2E, 0x3D, 0x3D, 0x2A, 0x3F, 0x4A, 0x5C, 0x23,
	0x11, 0x25, 0x2E, 0x00, 0x09, 0x27, 0x0A, 0x58, 0x34, 0x38, 0x3B, 0x5E,
	0x2F, 0x41, 0x18, 0x71, 0x3A, 0x15, 0x25, 0x1F, 0x36, 0x3B, 0x2D, 0x25,
	0x26, 0x1B, 0x35, 0x58, 0x59, 0x18, 0x0D, 0x3E, 0x58, 0x1E, 0x21, 0x77,
	0x22, 0x57, 0x19, 0x38, 0x38, 0x2D, 0x30, 0x57, 0x5B, 0x33, 0x36, 0x34,
	0x1C, 0x09, 0x32, 0x3A, 0x59, 0x23, 0x24, 0x74, 0x1D, 0x55, 0x21, 0x07,
	0x17, 0x1C, 0x39, 0x58, 0x0C, 0x1A, 0x3A, 0x39, 0x0C, 0x0A, 0x2B, 0x1A,
	0x3B, 0x22, 0x5C, 0x05, 0x1D, 0x26, 0x08, 0x13, 0x18, 0x22, 0x19, 0x59,
	0x20, 0x3A, 0x1B, 0x51, 0x00, 0x08, 0x06, 0x0F, 0x0F, 0x34, 0x19, 0x2B,
	0x59, 0x00, 0x08, 0x11, 0x74, 0x04, 0x0F, 0x0C, 0x44, 0x10, 0x02, 0x00,
	0x18, 0x18, 0x3A, 0x0D, 0x38, 0x0C, 0x39, 0x30, 0x0A, 0x4A, 0x5F, 0x5B,
	0x3A, 0x5E, 0x20, 0x17, 0x58, 0x05, 0x08, 0x0C, 0x22, 0x2E, 0x3B, 0x1C,
	0x17, 0x0F, 0x12, 0x18, 0x04, 0x33, 0x25, 0x08, 0x0E, 0x25, 0x28, 0x5B,
	0x33, 0x16, 0x27, 0x2D, 0x19, 0x22, 0x16, 0x2B, 0x53, 0x39, 0x0E, 0x11,
	0x0B, 0x57, 0x0A, 0x25, 0x0E, 0x5C, 0x39, 0x00, 0x0D, 0x36, 0x26, 0x59,
	0x38, 0x2E, 0x3A, 0x16, 0x58, 0x0A, 0x20, 0x7A, 0x0F, 0x23, 0x3E, 0x13,
	0x09, 0x00, 0x34, 0x29, 0x20, 0x73, 0x3B, 0x1B, 0x3C, 0x2C, 0x3B, 0x15,
	0x52, 0x29, 0x58, 0x0A, 0x3F, 0x52, 0x0B, 0x0A, 0x27, 0x0F, 0x26, 0x01,
	0x20, 0x0A, 0x36, 0x22, 0x0D, 0x38, 0x0E, 0x55, 0x18, 0x01, 0x5E, 0x17,
	0x02, 0x17, 0x3D, 0x5A, 0x77, 0x07, 0x50, 0x38, 0x1D, 0x01, 0x03, 0x53,
	0x02, 0x3D, 0x2B, 0x00, 0x2B, 0x00, 0x0E, 0x18, 0x04, 0x54, 0x3E, 0x21,
	0x0E, 0x5C, 0x06, 0x5C, 0x23, 0x76, 0x03, 0x23, 0x24, 0x33, 0x27, 0x1C,
	0x3B, 0x1E, 0x5D, 0x0F, 0x00, 0x05, 0x09, 0x31, 0x28, 0x1C, 0x11, 0x23,
	0x5A, 0x25, 0x3E, 0x29, 0x03, 0x21, 0x01, 0x5A, 0x05, 0x0F, 0x28, 0x15,
	0x19, 0x54, 0x18, 0x0F, 0x6D, 0x27, 0x4E, 0x5D, 0x3F, 0x0B, 0x03, 0x02,
	0x5B, 0x03, 0x07, 0x3B, 0x13, 0x3B, 0x58, 0x01, 0x0F, 0x0D, 0x34, 0x2E,
	0x16, 0x3D, 0x05, 0x34, 0x5D, 0x10, 0x0E, 0x12, 0x1E, 0x25, 0x31, 0x05,
	0x4A, 0x57, 0x5B, 0x73, 0x08, 0x39, 0x38, 0x09, 0x20, 0x55, 0x0F, 0x0B,
	0x12, 0x16, 0x1C, 0x2F, 0x0B, 0x58, 0x74, 0x15, 0x4E, 0x28, 0x2E, 0x1A,
	0x28, 0x50, 0x21, 0x1E, 0x06, 0x2F, 0x10, 0x57, 0x19, 0x76, 0x1F, 0x59,
	0x58, 0x09, 0x0E, 0x2B, 0x18, 0x0F, 0x0D, 0x2E, 0x5B, 0x20, 0x07, 0x5A,
	0x0A, 0x15, 0x0E, 0x1E, 0x2C, 0x69, 0x27, 0x26, 0x1D, 0x22, 0x2D, 0x54,
	0x38, 0x07, 0x1A, 0x0C, 0x5F, 0x12, 0x3C, 0x3A, 0x05, 0x3F, 0x0F, 0x07,
	0x06, 0x30, 0x5E, 0x03, 0x3B, 0x24, 0x17, 0x29, 0x26, 0x22, 0x3B, 0x03,
	0x28, 0x0A, 0x2C, 0x05, 0x3A, 0x38, 0x22, 0x1A, 0x29, 0x70, 0x04, 0x53,
	0x1C, 0x44, 0x09, 0x06, 0x08, 0x5C, 0x5B, 0x76, 0x25, 0x19, 0x03, 0x3F,
	0x74, 0x0D, 0x2A, 0x21, 0x59, 0x06, 0x5A, 0x0C, 0x5A, 0x38, 0x13, 0x0D,
	0x28, 0x26, 0x0A, 0x1A, 0x01, 0x29, 0x1E, 0x40, 0x71, 0x2E, 0x53, 0x05,
	0x08, 0x36, 0x3D, 0x50, 0x1D, 0x26, 0x0C, 0x22, 0x16, 0x3B, 0x29, 0x04,
	0x28, 0x34, 0x58, 0x11, 0x16, 0x0D, 0x33, 0x1D, 0x3E, 0x37, 0x5D, 0x2F,
	0x06, 0x23, 0x24, 0x5C, 0x0C, 0x01, 0x44, 0x32, 0x2A, 0x0C, 0x25, 0x11,
	0x33, 0x01, 0x52, 0x36, 0x31, 0x1A, 0x02, 0x4E, 0x34, 0x1A, 0x18, 0x2F,
	0x56, 0x3E, 0x20, 0x05, 0x06, 0x30, 0x04, 0x39, 0x36, 0x15, 0x2F, 0x5F,
	0x0D, 0x29, 0x15, 0x19, 0x3A, 0x5B, 0x75, 0x01, 0x31, 0x21, 0x21, 0x2C,
	0x1D, 0x4E, 0x3A, 0x5B, 0x0B, 0x05, 0x58, 0x26, 0x53, 0x1B, 0x55, 0x2B,
	0x05, 0x19, 0x0D, 0x38, 0x55, 0x1B, 0x1C, 0x37, 0x5C, 0x13, 0x18, 0x3D,
	0x11, 0x08, 0x11, 0x5F, 0x00, 0x73, 0x1C, 0x08, 0x14, 0x1B, 0x2F, 0x1B,
	0x53, 0x3A, 0x00, 0x2B, 0x1B, 0x15, 0x58, 0x03, 0x1B, 0x20, 0x2E, 0x41,
	0x1A, 0x33, 0x58, 0x2C, 0x2A, 0x3A, 0x73, 0x2F, 0x0A, 0x1A, 0x5B, 0x11,
	0x18, 0x00, 0x56, 0x40, 0x06, 0x03, 0x52, 0x01, 0x1C, 0x30, 0x04, 0x37,
	0x36, 0x0A, 0x35, 0x1F, 0x02, 0x2F, 0x02, 0x72, 0x04, 0x07, 0x39, 0x04,
	0x30, 0x35, 0x11, 0x07, 0x25, 0x0C, 0x23, 0x17, 0x17, 0x07, 0x27, 0x14,
	0x50, 0x0F, 0x2C, 0x0F, 0x23, 0x09, 0x09, 0x1A, 0x0D, 0x1B, 0x4A, 0x1F,
	0x3F, 0x0D, 0x35, 0x0A, 0x02, 0x3D, 0x34, 0x2A, 0x12, 0x5F, 0x3A, 0x69,
	0x0A, 0x18, 0x2D, 0x1F, 0x13, 0x2B, 0x31, 0x0A, 0x12, 0x0E, 0x5D, 0x54,
	0x14, 0x18, 0x1B, 0x39, 0x12, 0x5F, 0x26, 0x29, 0x38, 0x05, 0x01, 0x0E,
	0x75, 0x0A, 0x22, 0x58, 0x21, 0x0C, 0x08, 0x31, 0x26, 0x0C, 0x17, 0x16,
	0x59, 0x1A, 0x2E, 0x3A, 0x1A, 0x2D, 0x29, 0x23, 0x18, 0x07, 0x3B, 0x0C,
	0x3E, 0x15, 0x3C, 0x23, 0x1D, 0x2F, 0x1B, 0x5E, 0x50, 0x1D, 0x01, 0x18,
	0x21, 0x50, 0x3A, 0x1B, 0x73, 0x01, 0x13, 0x14, 0x00, 0x2D, 0x59, 0x15,
	0x24, 0x0F, 0x2C, 0x03, 0x00, 0x3C, 0x5C, 0x38, 0x05, 0x2F, 0x18, 0x20,
	0x73, 0x09, 0x19, 0x09, 0x0F, 0x11, 0x07, 0x2F, 0x45, 0x5C, 0x13, 0x5B,
	0x10, 0x1A, 0x2C, 0x13, 0x18, 0x05, 0x07, 0x02, 0x7A, 0x15, 0x10, 0x20,
	0x5A, 0x27, 0x5B, 0x14, 0x3A, 0x13, 0x13, 0x0E, 0x59, 0x0B, 0x0C, 0x69,
	0x0E, 0x28, 0x25, 0x28, 0x37, 0x5B, 0x56, 0x21, 0x29, 0x71, 0x00, 0x11,
	0x1C, 0x3F, 0x08, 0x3F, 0x0C, 0x1E, 0x2F, 0x36, 0x34, 0x56, 0x37, 0x20,
	0x17, 0x3F, 0x51, 0x0A, 0x23, 0x37, 0x08, 0x35, 0x39, 0x19, 0x30, 0x28,
	0x23, 0x09, 0x58, 0x75, 0x25, 0x37, 0x3C, 0x12, 0x11, 0x18, 0x31, 0x39,
	0x26, 0x29, 0x0B, 0x56, 0x09, 0x5D, 0x76, 0x20, 0x38, 0x3A, 0x22, 0x10,
	0x04, 0x0D, 0x22, 0x19, 0x71, 0x2B, 0x54, 0x1A, 0x3F, 0x06, 0x0A, 0x4A,
	0x21, 0x5C, 0x1A, 0x3A, 0x19, 0x3D, 0x5F, 0x27, 0x20, 0x14, 0x01, 0x44,
	0x3B, 0x58, 0x14, 0x00, 0x31, 0x25, 0x3F, 0x2B, 0x5C, 0x44, 0x3B, 0x0F,
	0x09, 0x37, 0x13, 0x74, 0x2D, 0x2A, 0x23, 0x3C, 0x17, 0x5C, 0x59, 0x08,
	0x0F, 0x73, 0x06, 0x27, 0x37, 0x3E, 0x70, 0x5E, 0x0F, 0x34, 0x1B, 0x12,
	0x38, 0x2C, 0x5B, 0x18, 0x2F, 0x02, 0x28, 0x05, 0x25, 0x10, 0x07, 0x07,
	0x2A, 0x3D, 0x14, 0x3F, 0x36, 0x08, 0x02, 0x0D, 0x47, 0x13, 0x2D, 0x5C,
	0x34, 0x54, 0x19, 0x39, 0x3E, 0x09, 0x3B, 0x50, 0x3C, 0x04, 0x37, 0x14,
	0x02, 0x18, 0x1B, 0x0A, 0x34, 0x50, 0x1F, 0x3E, 0x3A, 0x24, 0x04, 0x39,
	0x18, 0x20, 0x2E, 0x2D, 0x1B, 0x1A, 0x6D, 0x3D, 0x2B, 0x24, 0x5E, 0x75,
	0x2D, 0x36, 0x08, 0x0E, 0x00, 0x55, 0x22, 0x16, 0x5E, 0x07, 0x22, 0x18,
	0x24, 0x06, 0x0B, 0x15, 0x1B, 0x2A, 0x58, 0x20, 0x3B, 0x4A, 0x5B, 0x58,
	0x77, 0x3E, 0x39, 0x25, 0x01, 0x07, 0x1B, 0x54, 0x06, 0x0F, 0x31, 0x5B,
	0x36, 0x56, 0x07, 0x33, 0x26, 0x50, 0x27, 0x27, 0x28, 0x5F, 0x3B, 0x59,
	0x06, 0x36, 0x3C, 0x24, 0x5B, 0x00, 0x37, 0x26, 0x22, 0x24, 0x40, 0x7B,
	0x3A, 0x54, 0x3E, 0x27, 0x3A, 0x5F, 0x07, 0x07, 0x29, 0x7A, 0x5E, 0x34,
	0x00, 0x31, 0x34, 0x2B, 0x09, 0x02, 0x24, 0x0A, 0x05, 0x58, 0x0B, 0x0A,
	0x15, 0x3E, 0x58, 0x59, 0x3F, 0x74, 0x5C, 0x2A, 0x19, 0x52, 0x2A, 0x0B,
	0x02, 0x25, 0x04, 0x06, 0x00, 0x2A, 0x39, 0x38, 0x77, 0x02, 0x04, 0x1E,
	0x0C, 0x05, 0x14, 0x36, 0x2B, 0x07, 0x37, 0x05, 0x0F, 0x27, 0x1F, 0x0C,
	0x0F, 0x0D, 0x5A, 0x5F, 0x2E, 0x2F, 0x25, 0x39, 0x39, 0x1B, 0x3F, 0x3B,
	0x34, 0x07, 0x18, 0x24, 0x52, 0x26, 0x23, 0x2D, 0x02, 0x0C, 0x17, 0x33,
	0x20, 0x27, 0x0F, 0x36, 0x02, 0x18, 0x23, 0x33, 0x45, 0x3C, 0x0B, 0x1D,
	0x25, 0x25, 0x18, 0x20, 0x06, 0x0D, 0x0C, 0x2E, 0x35, 0x15, 0x56, 0x01,
	0x2F, 0x7B, 0x1E, 0x11, 0x25, 0x5D, 0x0C, 0x2F, 0x08, 0x3B, 0x5A, 0x15,
	0x18, 0x22, 0x08, 0x09, 0x2F, 0x22, 0x0E, 0x04, 0x31, 0x1A, 0x43, 0x33,
	0x5D, 0x3B, 0x05, 0x3C, 0x14, 0x36, 0x18, 0x14, 0x23, 0x02, 0x0D, 0x59,
	0x06, 0x36, 0x02, 0x01, 0x18, 0x7B, 0x2A, 0x05, 0x3C, 0x28, 0x0F, 0x38,
	0x37, 0x3C, 0x08, 0x06, 0x3F, 0x20, 0x01, 0x29, 0x21, 0x25, 0x00, 0x3D,
	0x2C, 0x20, 0x26, 0x2C, 0x3B, 0x1E, 0x09, 0x35, 0x0E, 0x37, 0x59, 0x3A,
	0x5E, 0x0E, 0x3A, 0x0D, 0x2C, 0x07, 0x00, 0x3D, 0x29, 0x18, 0x14, 0x09,
	0x29, 0x40, 0x34, 0x3A, 0x12, 0x00, 0x31, 0x24, 0x1D, 0x12, 0x22, 0x3B,
	0x08, 0x5A, 0x0B, 0x20, 0x5C, 0x2C, 0x2A, 0x27, 0x1E, 0x53, 0x27, 0x28,
	0x53, 0x0A, 0x3E, 0x72, 0x26, 0x0C, 0x16, 0x1F, 0x29, 0x2E, 0x52, 0x0B,
	0x3E, 0x2A, 0x3C, 0x2A, 0x3E, 0x38, 0x11, 0x2E, 0x37, 0x20, 0x1D, 0x2A,
	0x23, 0x29, 0x59, 0x02, 0x77, 0x35, 0x3B, 0x5C, 0x33, 0x06, 0x3C, 0x2D,
	0x5D, 0x2C, 0x23, 0x3B, 0x33, 0x1F, 0x0E, 0x11, 0x59, 0x00, 0x06, 0x00,
	0x74, 0x02, 0x27, 0x17, 0x1B, 0x04, 0x3E, 0x37, 0x02, 0x5F, 0x35, 0x1E,
	0x15, 0x5F, 0x1F, 0x14, 0x09, 0x52, 0x38, 0x3D, 0x7B, 0x0F, 0x2C, 0x0F,
	0x21, 0x0F, 0x58, 0x26, 0x14, 0x38, 0x05, 0x08, 0x29, 0x25, 0x00, 0x75,
	0x2E, 0x55, 0x5C, 0x11, 0x09, 0x07, 0x53, 0x57, 0x0F, 0x15, 0x08, 0x4A,
	0x3D, 0x44, 0x12, 0x0E, 0x12, 0x5F, 0x26, 0x25, 0x07, 0x14, 0x06, 0x28,
	0x32, 0x29, 0x0E, 0x02, 0x2D, 0x27, 0x1B, 0x2E, 0x0C, 0x3C, 0x71, 0x3D,
	0x0E, 0x17, 0x0D, 0x06, 0x1C, 0x39, 0x00, 0x08, 0x23, 0x06, 0x0B, 0x58,
	0x29, 0x01, 0x38, 0x37, 0x5F, 0x31, 0x09, 0x22, 0x34, 0x2D, 0x20, 0x30,
	0x06, 0x50, 0x3D, 0x0E, 0x21, 0x55, 0x30, 0x3E, 0x5E, 0x70, 0x05, 0x3B,
	0x0D, 0x44, 0x0C, 0x3F, 0x0F, 0x5F, 0x06, 0x24, 0x36, 0x00, 0x27, 0x3C,
	0x71, 0x5E, 0x53, 0x29, 0x00, 0x74, 0x19, 0x0B, 0x5F, 0x2F, 0x00, 0x25,
	0x38, 0x57, 0x40, 0x33, 0x07, 0x2B, 0x06, 0x0F, 0x6D, 0x07, 0x18, 0x41,
	0x08, 0x73, 0x1C, 0x31, 0x14, 0x3F, 0x05, 0x1A, 0x2E, 0x58, 0x12, 0x26,
	0x19, 0x13, 0x03, 0x53, 0x1B, 0x03, 0x2B, 0x07, 0x1B, 0x72, 0x07, 0x31,
	0x02, 0x32, 0x77, 0x16, 0x39, 0x2B, 0x31, 0x14, 0x58, 0x04, 0x3F, 0x52,
	0x74, 0x27, 0x4E, 0x05, 0x09, 0x2E, 0x35, 0x51, 0x3C, 0x3D, 0x15, 0x0F,
	0x05, 0x3F, 0x18, 0x6D, 0x22, 0x2A, 0x19, 0x2F, 0x35, 0x15, 0x03, 0x14,
	0x1F, 0x0D, 0x03, 0x37, 0x02, 0x2D, 0x04, 0x59, 0x19, 0x2B, 0x1B, 0x08,
	0x5E, 0x12, 0x3C, 0x12, 0x37, 0x3D, 0x04, 0x1C, 0x1D, 0x2C, 0x1D, 0x06,
	0x23, 0x09, 0x11, 0x1B, 0x0D, 0x06, 0x3F, 0x15, 0x15, 0x1B, 0x07, 0x2D,
	0x20, 0x1C, 0x35, 0x04, 0x0E, 0x2F, 0x5D, 0x07, 0x2B, 0x06, 0x17, 0x1F,
	0x2C, 0x5B, 0x22, 0x31, 0x19, 0x22, 0x5A, 0x3A, 0x09, 0x08, 0x2E, 0x34,
	0x26, 0x77, 0x25, 0x54, 0x01, 0x22, 0x0D, 0x3A, 0x57, 0x24, 0x40, 0x26,
	0x3D, 0x22, 0x37, 0x2F, 0x15, 0x5C, 0x23, 0x06, 0x28, 0x35, 0x18, 0x0C,
	0x25, 0x3B, 0x24, 0x3C, 0x2C, 0x5C, 0x5F, 0x2B, 0x07, 0x53, 0x3B, 0x38,
	0x2E, 0x23, 0x50, 0x1B, 0x08, 0x01, 0x08, 0x00, 0x0F, 0x11, 0x08, 0x38,
	0x33, 0x57, 0x01, 0x3A, 0x16, 0x06, 0x39, 0x3C, 0x10, 0x21, 0x37, 0x2C,
	0x2E, 0x3B, 0x1C, 0x2B, 0x5F, 0x01, 0x18, 0x5D, 0x0A, 0x1F, 0x28, 0x36,
	0x08, 0x00, 0x57, 0x06, 0x3A, 0x03, 0x56, 0x5F, 0x3A, 0x2F, 0x0E, 0x31,
	0x5F, 0x24, 0x07, 0x3B, 0x0D, 0x37, 0x3D, 0x25, 0x5A, 0x56, 0x2A, 0x1B,
	0x73, 0x59, 0x39, 0x3B, 0x2C, 0x04, 0x1B, 0x18, 0x3B, 0x1D, 0x0A, 0x54,
	0x59, 0x14, 0x0C, 0x27, 0x14, 0x05, 0x3B, 0x0A, 0x37, 0x2A, 0x31, 0x20,
	0x1A, 0x20, 0x14, 0x0D, 0x5B, 0x0C, 0x09, 0x14, 0x18, 0x07, 0x40, 0x38,
	0x03, 0x54, 0x27, 0x5D, 0x2E, 0x0F, 0x28, 0x56, 0x3D, 0x11, 0x55, 0x3B,
	0x16, 0x3E, 0x27, 0x1A, 0x2C, 0x21, 0x0A, 0x1A, 0x23, 0x10, 0x34, 0x26,
	0x2F, 0x3F, 0x50, 0x5A, 0x2F, 0x33, 0x3E, 0x04, 0x00, 0x5B, 0x69, 0x28,
	0x20, 0x45, 0x0F, 0x71, 0x2A, 0x0E, 0x0A, 0x13, 0x10, 0x22, 0x51, 0x37,
	0x1F, 0x73, 0x5E, 0x05, 0x57, 0x0A, 0x37, 0x00, 0x0C, 0x0A, 0x03, 0x3B,
	0x07, 0x17, 0x59, 0x04, 0x69, 0x55, 0x00, 0x04, 0x09, 0x01, 0x09, 0x18,
	0x0D, 0x53, 0x04, 0x1D, 0x07, 0x3F, 0x1C, 0x05, 0x3A, 0x57, 0x38, 0x39,
	0x21, 0x5E, 0x37, 0x3D, 0x32, 0x2B, 0x0B, 0x56, 0x1F, 0x3F, 0x2F, 0x16,
	0x53, 0x22, 0x5D, 0x38, 0x0F, 0x2B, 0x59, 0x3E, 0x2D, 0x2A, 0x29, 0x5D,
	0x38, 0x2D, 0x2F, 0x03, 0x00, 0x11, 0x1A, 0x0D, 0x35, 0x1A, 0x53, 0x10,
	0x18, 0x27, 0x3D, 0x5C, 0x70, 0x1B, 0x55, 0x36, 0x5A, 0x74, 0x08, 0x0C,
	0x41, 0x53, 0x15, 0x19, 0x50, 0x0F, 0x3A, 0x2A, 0x2A, 0x26, 0x20, 0x2E,
	0x32, 0x2A, 0x54, 0x24, 0x26, 0x75, 0x3A, 0x13, 0x17, 0x29, 0x76, 0x1A,
	0x12, 0x1F, 0x52, 0x14, 0x3F, 0x4E, 0x5E, 0x1C, 0x31, 0x3A, 0x0B, 0x2B,
	0x0F, 0x1A, 0x19, 0x06, 0x5B, 0x22, 0x75, 0x08, 0x2D, 0x1D, 0x32, 0x0E,
	0x0A, 0x28, 0x38, 0x39, 0x36, 0x07, 0x00, 0x5A, 0x13, 0x76, 0x21, 0x0A,
	0x03, 0x53, 0x3B, 0x55, 0x00, 0x05, 0x21, 0x70, 0x58, 0x55, 0x41, 0x38,
	0x23, 0x2B, 0x38, 0x04, 0x19, 0x2D, 0x07, 0x0E, 0x03, 0x3A, 0x10, 0x05,
	0x27, 0x3D, 0x12, 0x13, 0x27, 0x07, 0x1F, 0x0F, 0x34, 0x5F, 0x33, 0x1F,
	0x02, 0x28, 0x00, 0x2E, 0x0A, 0x04, 0x27, 0x54, 0x2D, 0x1D, 0x59, 0x36,
	0x20, 0x11, 0x09, 0x3E, 0x14, 0x24, 0x20, 0x3A, 0x31, 0x15, 0x15, 0x54,
	0x0D, 0x12, 0x7B, 0x36, 0x35, 0x3F, 0x39, 0x09, 0x02, 0x32, 0x2C, 0x3C,
	0x31, 0x14, 0x27, 0x38, 0x25, 0x2C, 0x19, 0x3B, 0x3D, 0x5A, 0x2E, 0x1C,
	0x2E, 0x05, 0x3C, 0x20, 0x5C, 0x26, 0x5B, 0x59, 0x26, 0x1D, 0x30, 0x2C,
	0x18, 0x03, 0x25, 0x0F, 0x2A, 0x05, 0x2F, 0x1E, 0x55, 0x0A, 0x04, 0x15,
	0x5A, 0x0B, 0x0F, 0x06, 0x14, 0x0F, 0x16, 0x18, 0x1A, 0x74, 0x29, 0x0B,
	0x2F, 0x5D, 0x0D, 0x08, 0x4E, 0x0B, 0x2E, 0x15, 0x58, 0x35, 0x23, 0x3F,
	0x2B, 0x09, 0x52, 0x3E, 0x18, 0x70, 0x0A, 0x57, 0x45, 0x1C, 0x01, 0x15,
	0x13, 0x04, 0x28, 0x2B, 0x18, 0x59, 0x2C, 0x39, 0x7B, 0x1F, 0x08, 0x03,
	0x2D, 0x6D, 0x0E, 0x0B, 0x2C, 0x06, 0x23, 0x59, 0x2A, 0x19, 0x2A, 0x0F,
	0x34, 0x34, 0x5A, 0x26, 0x31, 0x26, 0x12, 0x5F, 0x18, 0x28, 0x27, 0x03,
	0x16, 0x3E, 0x33, 0x5B, 0x12, 0x18, 0x0D, 0x14, 0x3F, 0x25, 0x0B, 0x1D,
	0x31, 0x23, 0x0F, 0x03, 0x44, 0x7B, 0x0B, 0x0E, 0x3A, 0x5C, 0x08, 0x06,
	0x18, 0x24, 0x3F, 0x36, 0x15, 0x2C, 0x1E, 0x28, 0x7B, 0x2F, 0x38, 0x2B,
	0x25, 0x29, 0x05, 0x34, 0x39, 0x5E, 0x38, 0x21, 0x06, 0x0D, 0x59, 0x11,
	0x0F, 0x57, 0x0C, 0x31, 0x27, 0x0D, 0x52, 0x1E, 0x29, 0x31, 0x59, 0x4A,
	0x3F, 0x21, 0x34, 0x29, 0x35, 0x5F, 0x5A, 0x00, 0x47, 0x4E, 0x41, 0x21,
	0x38, 0x05, 0x58, 0x1A, 0x2E, 0x25, 0x0A, 0x27, 0x20, 0x05, 0x14, 0x5B,
	0x15, 0x36, 0x1D, 0x0A, 0x05, 0x30, 0x06, 0x32, 0x7B, 0x3B, 0x4A, 0x22,
	0x3A, 0x1B, 0x47, 0x34, 0x58, 0x5B, 0x10, 0x01, 0x37, 0x58, 0x25, 0x14,
	0x38, 0x15, 0x25, 0x1A, 0x3A, 0x3F, 0x3B, 0x1D, 0x3B, 0x30, 0x01, 0x53,
	0x5B, 0x0E, 0x6D, 0x27, 0x35, 0x45, 0x13, 0x30, 0x47, 0x56, 0x0C, 0x3F,
	0x0B, 0x0F, 0x08, 0x5F, 0x44, 0x6D, 0x04, 0x55, 0x16, 0x0E, 0x33, 0x1B,
	0x02, 0x01, 0x59, 0x11, 0x14, 0x2D, 0x03, 0x32, 0x2D, 0x28, 0x20, 0x1A,
	0x0E, 0x31, 0x3E, 0x2B, 0x27, 0x04, 0x2F, 0x00, 0x26, 0x0C, 0x00, 0x2E,
	0x07, 0x04, 0x26, 0x2A, 0x28, 0x1F, 0x57, 0x02, 0x28, 0x77, 0x5C, 0x24,
	0x3C, 0x3D, 0x0C, 0x35, 0x32, 0x02, 0x0E, 0x7B, 0x54, 0x57, 0x0A, 0x1A,
	0x34, 0x3B, 0x31, 0x36, 0x39, 0x2C, 0x05, 0x2F, 0x2F, 0x31, 0x30, 0x07,
	0x06, 0x36, 0x3B, 0x12, 0x39, 0x4A, 0x41, 0x32, 0x70, 0x07, 0x09, 0x57,
	0x0A, 0x23, 0x5D, 0x35, 0x0B, 0x09, 0x69, 0x28, 0x08, 0x3B, 0x5C, 0x3A,
	0x2A, 0x14, 0x02, 0x3E, 0x6D, 0x01, 0x2E, 0x0F, 0x28, 0x23, 0x2F, 0x2D,
	0x07, 0x19, 0x2B, 0x1E, 0x53, 0x36, 0x2E, 0x32, 0x15, 0x38, 0x22, 0x19,
	0x31, 0x2B, 0x00, 0x3C, 0x21, 0x34, 0x05, 0x2E, 0x3B, 0x26, 0x13, 0x5E,
	0x34, 0x0C, 0x01, 0x09, 0x38, 0x1B, 0x0D, 0x27, 0x24, 0x36, 0x19, 0x22,
	0x00, 0x70, 0x14, 0x3B, 0x14, 0x27, 0x28, 0x5A, 0x25, 0x28, 0x1C, 0x23,
	0x21, 0x13, 0x38, 0x2D, 0x18, 0x21, 0x55, 0x3C, 0x5C, 0x2A, 0x1A, 0x2A,
	0x25, 0x1F, 0x33, 0x0E, 0x2B, 0x28, 0x2D, 0x29, 0x1E, 0x11, 0x29, 0x27,
	0x0C, 0x25, 0x13, 0x05, 0x31, 0x28, 0x0E, 0x35, 0x3C, 0x40, 0x0F, 0x06,
	0x18, 0x37, 0x1A, 0x33, 0x2A, 0x2D, 0x08, 0x25, 0x72, 0x25, 0x0D, 0x5E,
	0x5C, 0x1B, 0x34, 0x0A, 0x25, 0x0C, 0x12, 0x2A, 0x32, 0x21, 0x13, 0x01,
	0x3F, 0x57, 0x08, 0x3A, 0x08, 0x25, 0x11, 0x20, 0x3E, 0x73, 0x39, 0x34,
	0x2A, 0x3D, 0x04, 0x0A, 0x27, 0x39, 0x3C, 0x08, 0x2F, 0x55, 0x18, 0x0A,
	0x71, 0x23, 0x07, 0x3B, 0x3A, 0x30, 0x38, 0x05, 0x36, 0x3E, 0x2D, 0x1B,
	0x03, 0x14, 0x3A, 0x24, 0x18, 0x32, 0x0F, 0x39, 0x31, 0x54, 0x2E, 0x23,
	0x52, 0x0B, 0x16, 0x53, 0x2F, 0x5C, 0x71, 0x1F, 0x29, 0x00, 0x3D, 0x21,
	0x3B, 0x30, 0x29, 0x3C, 0x05, 0x3C, 0x16, 0x3F, 0x1B, 0x23, 0x1A, 0x39,
	0x0C, 0x2D, 0x09, 0x47, 0x10, 0x03, 0x2E, 0x29, 0x09, 0x10, 0x06, 0x20,
	0x73, 0x5B, 0x2D, 0x1E, 0x18, 0x31, 0x01, 0x0B, 0x28, 0x5D, 0x37, 0x14,
	0x2D, 0x1D, 0x01, 0x2D, 0x01, 0x37, 0x36, 0x1B, 0x13, 0x3A, 0x4A, 0x24,
	0x23, 0x77, 0x35, 0x33, 0x2B, 0x13, 0x23, 0x2A, 0x20, 0x0F, 0x5B, 0x08,
	0x01, 0x0C, 0x16, 0x3F, 0x05, 0x18, 0x0D, 0x5B, 0x5F, 0x01, 0x2B, 0x0A,
	0x26, 0x3C, 0x09, 0x55, 0x50, 0x57, 0x1F, 0x29, 0x19, 0x58, 0x18, 0x0A,
	0x06, 0x5F, 0x13, 0x58, 0x3E, 0x14, 0x01, 0x28, 0x27, 0x0C, 0x33, 0x3F,
	0x03, 0x26, 0x52, 0x16, 0x29, 0x50, 0x5F, 0x5D, 0x25, 0x24, 0x13, 0x26,
	0x38, 0x2C, 0x5C, 0x57, 0x2F, 0x20, 0x13, 0x5D, 0x34, 0x28, 0x31, 0x00,
	0x07, 0x34, 0x58, 0x1B, 0x32, 0x5E, 0x16, 0x03, 0x3D, 0x7B, 0x21, 0x57,
	0x08, 0x29, 0x72, 0x20, 0x30, 0x34, 0x1E, 0x1A, 0x16, 0x25, 0x1A, 0x38,
	0x69, 0x09, 0x1B, 0x0D, 0x21, 0x07, 0x1B, 0x4E, 0x3B, 0x03, 0x1A, 0x35,
	0x38, 0x23, 0x01, 0x15, 0x16, 0x1B, 0x23, 0x06, 0x03, 0x19, 0x58, 0x06,
	0x18, 0x30, 0x29, 0x34, 0x5D, 0x19, 0x2F, 0x38, 0x19, 0x2D, 0x06, 0x23,
	0x35, 0x13, 0x21, 0x1F, 0x09, 0x36, 0x32, 0x3F, 0x29, 0x30, 0x3E, 0x32,
	0x1A, 0x3C, 0x37, 0x2F, 0x36, 0x1F, 0x24, 0x69, 0x0F, 0x1B, 0x34, 0x0F,
	0x17, 0x19, 0x10, 0x45, 0x18, 0x29, 0x02, 0x0D, 0x20, 0x0E, 0x14, 0x18,
	0x2E, 0x2D, 0x3D, 0x09, 0x2A, 0x33, 0x29, 0x59, 0x34, 0x1A, 0x0D, 0x2F,
	0x18, 0x33, 0x15, 0x08, 0x2C, 0x1A, 0x0F, 0x1D, 0x59, 0x04, 0x5A, 0x38,
	0x5D, 0x08, 0x07, 0x52, 0x70, 0x15, 0x0C, 0x0F, 0x04, 0x2C, 0x27, 0x0A,
	0x2D, 0x03, 0x15, 0x55, 0x22, 0x14, 0x13, 0x0D, 0x0B, 0x0A, 0x5B, 0x1A,
	0x16, 0x5C, 0x04, 0x58, 0x1A, 0x2B, 0x0A, 0x39, 0x57, 0x21, 0x08, 0x0F,
	0x13, 0x1C, 0x29, 0x23, 0x5D, 0x0D, 0x26, 0x3B, 0x31, 0x07, 0x0C, 0x17,
	0x5F, 0x0D, 0x38, 0x00, 0x17, 0x20, 0x13, 0x09, 0x22, 0x27, 0x3B, 0x04,
	0x0A, 0x2A, 0x20, 0x2C, 0x71, 0x3B, 0x54, 0x5B, 0x3F, 0x0A, 0x22, 0x33,
	0x0B, 0x23, 0x27, 0x06, 0x2D, 0x24, 0x0F, 0x15, 0x22, 0x19, 0x3B, 0x01,
	0x05, 0x07, 0x2C, 0x34, 0x40, 0x76, 0x3D, 0x54, 0x5B, 0x06, 0x29, 0x55,
	0x05, 0x0B, 0x24, 0x1B, 0x01, 0x14, 0x16, 0x58, 0x36, 0x1A, 0x39, 0x20,
	0x33, 0x25, 0x23, 0x0F, 0x0A, 0x29, 0x0A, 0x3C, 0x02, 0x23, 0x22, 0x3B,
	0x3A, 0x0F, 0x58, 0x11, 0x05, 0x16, 0x39, 0x3C, 0x1B, 0x14, 0x04, 0x24,
	0x08, 0x38, 0x28, 0x09, 0x57, 0x5E, 0x2A, 0x16, 0x0E, 0x0D, 0x00, 0x19,
	0x10, 0x18, 0x14, 0x28, 0x3F, 0x05, 0x5C, 0x52, 0x56, 0x5A, 0x70, 0x5C,
	0x2D, 0x5B, 0x3C, 0x3A, 0x3B, 0x12, 0x2A, 0x1B, 0x11, 0x25, 0x51, 0x06,
	0x18, 0x25, 0x35, 0x00, 0x5F, 0x33, 0x23, 0x3F, 0x11, 0x3C, 0x3A, 0x0F,
	0x5A, 0x3B, 0x1E, 0x0E, 0x00, 0x3A, 0x0F, 0x5E, 0x3C, 0x33, 0x5A, 0x35,
	0x21, 0x2E, 0x36, 0x0B, 0x26, 0x3F, 0x1A, 0x24, 0x0A, 0x2E, 0x28, 0x12,
	0x74, 0x27, 0x56, 0x5D, 0x31, 0x34, 0x09, 0x16, 0x34, 0x2A, 0x0D, 0x0F,
	0x12, 0x41, 0x58, 0x0C, 0x05, 0x32, 0x1E, 0x09, 0x2A, 0x25, 0x3B, 0x0F,
	0x1E, 0x37, 0x34, 0x2C, 0x04, 0x39, 0x37, 0x01, 0x33, 0x17, 0x53, 0x30,
	0x26, 0x18, 0x18, 0x20, 0x06, 0x07, 0x59, 0x05, 0x0F, 0x74, 0x2F, 0x2F,
	0x34, 0x05, 0x0C, 0x3E, 0x03, 0x36, 0x31, 0x38, 0x34, 0x57, 0x25, 0x0E,
	0x07, 0x03, 0x0C, 0x21, 0x12, 0x37, 0x43, 0x33, 0x0A, 0x2F, 0x2F, 0x19,
	0x19, 0x57, 0x1C, 0x25, 0x5B, 0x00, 0x1F, 0x1A, 0x01, 0x29, 0x26, 0x0A,
	0x02, 0x70, 0x16, 0x35, 0x25, 0x0A, 0x13, 0x5B, 0x29, 0x29, 0x5D, 0x23,
	0x58, 0x58, 0x21, 0x1F, 0x17, 0x59, 0x23, 0x5B, 0x3B, 0x2C, 0x19, 0x32,
	0x0D, 0x40, 0x05, 0x47, 0x39, 0x2A, 0x3B, 0x04, 0x01, 0x11, 0x18, 0x3C,
	0x08, 0x0A, 0x00, 0x3D, 0x19, 0x33, 0x39, 0x15, 0x0A, 0x26, 0x26, 0x5D,
	0x18, 0x36, 0x0A, 0x73, 0x5C, 0x06, 0x5E, 0x1A, 0x73, 0x54, 0x18, 0x3E,
	0x24, 0x06, 0x24, 0x09, 0x17, 0x01, 0x03, 0x19, 0x59, 0x1B, 0x11, 0x34,
	0x1C, 0x06, 0x21, 0x07, 0x2B, 0x36, 0x0D, 0x16, 0x22, 0x38, 0x25, 0x54,
	0x1A, 0x04, 0x76, 0x2B, 0x00, 0x1D, 0x3C, 0x7A, 0x2F, 0x37, 0x0F, 0x3D,
	0x2F, 0x05, 0x18, 0x0F, 0x24, 0x32, 0x23, 0x27, 0x1C, 0x2D, 0x01, 0x05,
	0x0B, 0x36, 0x26, 0x2E, 0x08, 0x35, 0x25, 0x26, 0x13, 0x59, 0x27, 0x45,
	0x39, 0x33, 0x5E, 0x00, 0x0B, 0x52, 0x14, 0x01, 0x19, 0x00, 0x5D, 0x2E,
	0x08, 0x0D, 0x39, 0x3A, 0x72, 0x47, 0x56, 0x3A, 0x25, 0x16, 0x1C, 0x2E,
	0x5F, 0x31, 0x35, 0x36, 0x53, 0x0B, 0x53, 0x14, 0x02, 0x0D, 0x07, 0x5C,
	0x28, 0x58, 0x4A, 0x2A, 0x12, 0x0C, 0x14, 0x0C, 0x07, 0x25, 0x14, 0x0A,
	0x0A, 0x1B, 0x13, 0x7B, 0x03, 0x52, 0x41, 0x07, 0x21, 0x38, 0x2F, 0x1E,
	0x1C, 0x32, 0x5C, 0x35, 0x39, 0x05, 0x06, 0x01, 0x33, 0x1C, 0x2E, 0x32,
	0x5D, 0x06, 0x17, 0x24, 0x72, 0x09, 0x50, 0x09, 0x32, 0x35, 0x26, 0x56,
	0x1F, 0x0E, 0x34, 0x47, 0x54, 0x18, 0x40, 0x72, 0x5D, 0x2B, 0x58, 0x1B,
	0x0D, 0x39, 0x03, 0x1F, 0x1C, 0x10, 0x14, 0x0F, 0x03, 0x38, 0x35, 0x24,
	0x19, 0x58, 0x07, 0x32, 0x59, 0x2E, 0x16, 0x1B, 0x20, 0x14, 0x00, 0x17,
	0x5D, 0x35, 0x47, 0x31, 0x36, 0x22, 0x36, 0x29, 0x1B, 0x5C, 0x2C, 0x0D,
	0x14, 0x3B, 0x3C, 0x3C, 0x0A, 0x5D, 0x30, 0x2C, 0x13, 0x26, 0x3E, 0x59,
	0x23, 0x26, 0x32, 0x28, 0x58, 0x41, 0x38, 0x31, 0x5B, 0x37, 0x34, 0x24,
	0x32, 0x35, 0x23, 0x34, 0x44, 0x2D, 0x0A, 0x39, 0x16, 0x38, 0x28, 0x38,
	0x4A, 0x01, 0x29, 0x00, 0x04, 0x56, 0x00, 0x3B, 0x15, 0x35, 0x23, 0x39,
	0x03, 0x71, 0x25, 0x2A, 0x0A, 0x02, 0x7B, 0x04, 0x33, 0x1F, 0x33, 0x0E,
	0x36, 0x2A, 0x38, 0x33, 0x74, 0x1F, 0x08, 0x20, 0x3E, 0x30, 0x22, 0x09,
	0x3A, 0x3E, 0x14, 0x1F, 0x2E, 0x06, 0x5E, 0x0E, 0x02, 0x2B, 0x06, 0x01,
	0x1A, 0x0B, 0x0A, 0x2D, 0x3E, 0x38, 0x09, 0x2B, 0x36, 0x5F, 0x72, 0x0A,
	0x13, 0x5E, 0x1A, 0x1A, 0x2E, 0x58, 0x36, 0x0C, 0x0F, 0x3F, 0x15, 0x07,
	0x1E, 0x31, 0x0B, 0x53, 0x0F, 0x21, 0x34, 0x01, 0x04, 0x0A, 0x33, 0x32,
	0x0F, 0x2D, 0x22, 0x09, 0x71, 0x2A, 0x0E, 0x1A, 0x04, 0x38, 0x0A, 0x12,
	0x0C, 0x53, 0x13, 0x22, 0x15, 0x39, 0x2C, 0x0F, 0x3E, 0x53, 0x09, 0x5B,
	0x1A, 0x24, 0x2F, 0x17, 0x5A, 0x70, 0x3B, 0x02, 0x19, 0x53, 0x23, 0x28,
	0x09, 0x1C, 0x33, 0x6D, 0x5E, 0x15, 0x1B, 0x22, 0x37, 0x0F, 0x3B, 0x1D,
	0x1B, 0x36, 0x5C, 0x04, 0x0C, 0x3C, 0x10, 0x34, 0x2F, 0x0C, 0x2E, 0x0F,
	0x5B, 0x03, 0x1F, 0x08, 0x0F, 0x0A, 0x34, 0x1F, 0x52, 0x24, 0x36, 0x0C,
	0x57, 0x09, 0x16, 0x19, 0x56, 0x58, 0x1C, 0x0D, 0x5B, 0x03, 0x17, 0x00,
	0x26, 0x26, 0x57, 0x1E, 0x02, 0x0D, 0x26, 0x58, 0x3F, 0x13, 0x2A, 0x03,
	0x32, 0x3C, 0x5B, 0x0F, 0x59, 0x55, 0x17, 0x2E, 0x28, 0x0B, 0x57, 0x0A,
	0x3C, 0x69, 0x43, 0x34, 0x07, 0x32, 0x34, 0x3A, 0x00, 0x1B, 0x07, 0x2B,
	0x09, 0x11, 0x41, 0x32, 0x38, 0x26, 0x23, 0x29, 0x58, 0x16, 0x25, 0x13,
	0x29, 0x02, 0x11, 0x59, 0x29, 0x14, 0x29, 0x71, 0x23, 0x37, 0x0F, 0x1F,
	0x71, 0x1C, 0x28, 0x5A, 0x3A, 0x37, 0x25, 0x4E, 0x59, 0x2C, 0x04, 0x5C,
	0x15, 0x1E, 0x59, 0x29, 0x1E, 0x0F, 0x25, 0x11, 0x15, 0x0D, 0x0D, 0x36,
	0x13, 0x08, 0x09, 0x19, 0x20, 0x11, 0x77, 0x2F, 0x58, 0x2B, 0x1B, 0x0C,
	0x55, 0x58, 0x37, 0x06, 0x14, 0x36, 0x26, 0x0A, 0x21, 0x03, 0x20, 0x0B,
	0x24, 0x24, 0x35, 0x00, 0x03, 0x1C, 0x52, 0x09, 0x1F, 0x0D, 0x0A, 0x27,
	0x69, 0x5D, 0x0F, 0x38, 0x33, 0x26, 0x03, 0x57, 0x29, 0x38, 0x27, 0x07,
	0x03, 0x1A, 0x39, 0x0F, 0x0F, 0x58, 0x39, 0x1B, 0x03, 0x14, 0x12, 0x04,
	0x2C, 0x3A, 0x26, 0x59, 0x05, 0x5D, 0x17, 0x38, 0x12, 0x29, 0x24, 0x21,
	0x23, 0x02, 0x23, 0x1F, 0x16, 0x2B, 0x37, 0x03, 0x3B, 0x75, 0x03, 0x50,
	0x45, 0x00, 0x69, 0x15, 0x13, 0x1F, 0x2E, 0x7B, 0x34, 0x56, 0x29, 0x31,
	0x15, 0x1C, 0x12, 0x08, 0x31, 0x0A, 0x08, 0x02, 0x01, 0x12, 0x0E, 0x21,
	0x0B, 0x09, 0x59, 0x75, 0x5D, 0x24, 0x3A, 0x2D, 0x34, 0x0A, 0x37, 0x3A,
	0x31, 0x24, 0x09, 0x03, 0x2B, 0x38, 0x2E, 0x1E, 0x53, 0x5D, 0x3B, 0x0A,
	0x54, 0x53, 0x1F, 0x07, 0x74, 0x5A, 0x2C, 0x21, 0x05, 0x10, 0x1B, 0x10,
	0x3A, 0x59, 0x27, 0x0E, 0x57, 0x3B, 0x33, 0x0A, 0x35, 0x2C, 0x14, 0x2E,
	0x30, 0x39, 0x50, 0x3B, 0x0F, 0x26, 0x27, 0x28, 0x5C, 0x3E, 0x3B, 0x05,
	0x1B, 0x58, 0x20, 0x00, 0x3E, 0x50, 0x0A, 0x27, 0x38, 0x07, 0x37, 0x00,
	0x0E, 0x76, 0x04, 0x07, 0x3E, 0x38, 0x74, 0x5D, 0x03, 0x1F, 0x1C, 0x70,
	0x38, 0x54, 0x5F, 0x1C, 0x15, 0x2D, 0x05, 0x06, 0x09, 0x11, 0x25, 0x32,
	0x24, 0x1A, 0x72, 0x22, 0x28, 0x04, 0x24, 0x07, 0x36, 0x38, 0x5E, 0x2E,
	0x0F, 0x55, 0x53, 0x1E, 0x32, 0x3A, 0x5A, 0x36, 0x0B, 0x25, 0x36, 0x0A,
	0x0A, 0x5D, 0x3F, 0x72, 0x29, 0x02, 0x34, 0x39, 0x31, 0x0B, 0x33, 0x1F,
	0x53, 0x28, 0x1E, 0x02, 0x24, 0x23, 0x05, 0x0E, 0x03, 0x34, 0x5B, 0x29,
	0x38, 0x06, 0x3C, 0x13, 0x31, 0x1E, 0x08, 0x38, 0x1E, 0x24, 0x2E, 0x0C,
	0x14, 0x2C, 0x2D, 0x02, 0x4A, 0x5F, 0x1B, 0x31, 0x0A, 0x2E, 0x36, 0x28,
	0x27, 0x21, 0x0C, 0x57, 0x52, 0x01, 0x0F, 0x27, 0x2F, 0x40, 0x11, 0x01,
	0x04, 0x58, 0x2D, 0x7B, 0x5E, 0x0D, 0x38, 0x09, 0x71, 0x5A, 0x17, 0x1A,
	0x21, 0x0F, 0x1C, 0x52, 0x3E, 0x05, 0x16, 0x28, 0x25, 0x2F, 0x32, 0x75,
	0x34, 0x51, 0x36, 0x5F, 0x75, 0x06, 0x26, 0x41, 0x3E, 0x0F, 0x59, 0x00,
	0x39, 0x0D, 0x07, 0x2D, 0x2C, 0x5A, 0x2C, 0x76, 0x3A, 0x35, 0x41, 0x3D,
	0x29, 0x28, 0x1B, 0x3E, 0x0A, 0x04, 0x08, 0x10, 0x1A, 0x0A, 0x31, 0x07,
	0x2E, 0x27, 0x5D, 0x0D, 0x14, 0x08, 0x0C, 0x40, 0x0C, 0x43, 0x2D, 0x5C,
	0x26, 0x76, 0x59, 0x03, 0x1F, 0x1B, 0x01, 0x3F, 0x2A, 0x36, 0x11, 0x34,
	0x26, 0x12, 0x29, 0x1A, 0x36, 0x3F, 0x50, 0x06, 0x1F, 0x70, 0x16, 0x08,
	0x2A, 0x1E, 0x31, 0x07, 0x25, 0x3A, 0x01, 0x2E, 0x26, 0x56, 0x27, 0x1A,
	0x2F, 0x47, 0x14, 0x1F, 0x0E, 0x00, 0x2A, 0x59, 0x36, 0x44, 0x18, 0x2E,
	0x12, 0x29, 0x1A, 0x06, 0x5A, 0x30, 0x1C, 0x40, 0x34, 0x07, 0x2E, 0x18,
	0x3F, 0x05, 0x3F, 0x0F, 0x2C, 0x2A, 0x00, 0x35, 0x0E, 0x0A, 0x3F, 0x37,
	0x34, 0x53, 0x0D, 0x5A, 0x74, 0x01, 0x50, 0x0C, 0x5F, 0x38, 0x1C, 0x17,
	0x45, 0x04, 0x14, 0x1C, 0x3B, 0x14, 0x59, 0x18, 0x14, 0x59, 0x36, 0x2A,
	0x72, 0x3C, 0x37, 0x17, 0x58, 0x15, 0x3F, 0x19, 0x1A, 0x28, 0x74, 0x0D,
	0x34, 0x5B, 0x2C, 0x0B, 0x47, 0x26, 0x1A, 0x02, 0x3B, 0x58, 0x23, 0x0D,
	0x04, 0x14, 0x22, 0x2E, 0x16, 0x2C, 0x00, 0x06, 0x38, 0x5B, 0x02, 0x0D,
	0x29, 0x35, 0x06, 0x28, 0x2B, 0x2F, 0x17, 0x23, 0x5D, 0x10, 0x5D, 0x35,
	0x29, 0x0F, 0x15, 0x2B, 0x15, 0x3C, 0x3D, 0x1B, 0x39, 0x52, 0x5D, 0x3A,
	0x21, 0x5F, 0x23, 0x20, 0x18, 0x30, 0x3E, 0x3B, 0x16, 0x18, 0x7B, 0x21,
	0x3B, 0x14, 0x2E, 0x38, 0x00, 0x50, 0x00, 0x0D, 0x07, 0x06, 0x36, 0x38,
	0x24, 0x2F, 0x3F, 0x23, 0x24, 0x2D, 0x37, 0x35, 0x2E, 0x22, 0x21, 0x04,
	0x5C, 0x16, 0x14, 0x06, 0x74, 0x0D, 0x07, 0x25, 0x24, 0x7B, 0x2B, 0x0A,
	0x16, 0x1E, 0x26, 0x0E, 0x0C, 0x28, 0x3C, 0x16, 0x43, 0x15, 0x2B, 0x08,
	0x37, 0x06, 0x15, 0x17, 0x0A, 0x30, 0x39, 0x2B, 0x56, 0x2D, 0x09, 0x5F,
	0x15, 0x3A, 0x33, 0x76, 0x5E, 0x2D, 0x2C, 0x5A, 0x36, 0x02, 0x0F, 0x0F,
	0x3C, 0x11, 0x36, 0x2F, 0x0D, 0x12, 0x1A, 0x5F, 0x2C, 0x07, 0x5C, 0x05,
	0x0D, 0x3B, 0x0F, 0x52, 0x15, 0x58, 0x28, 0x04, 0x1E, 0x3B, 0x5A, 0x34,
	0x3E, 0x1A, 0x0B, 0x3C, 0x1B, 0x5A, 0x3A, 0x10, 0x19, 0x57, 0x00, 0x27,
	0x36, 0x3E, 0x13, 0x23, 0x0A, 0x27, 0x1E, 0x14, 0x2C, 0x03, 0x2D, 0x5D,
	0x17, 0x0A, 0x05, 0x06, 0x54, 0x03, 0x26, 0x5B, 0x06, 0x03, 0x0D, 0x21,
	0x1E, 0x15, 0x19, 0x33, 0x1C, 0x3E, 0x0A, 0x3A, 0x03, 0x16, 0x5F, 0x35,
	0x1C, 0x13, 0x26, 0x22, 0x29, 0x0E, 0x0C, 0x1D, 0x38, 0x2A, 0x2A, 0x53,
	0x1E, 0x5C, 0x36, 0x36, 0x19, 0x00, 0x32, 0x06, 0x35, 0x14, 0x00, 0x40,
	0x10, 0x54, 0x07, 0x07, 0x53, 0x1A, 0x23, 0x2D, 0x14, 0x3C, 0x18, 0x09,
	0x51, 0x3A, 0x2F, 0x14, 0x5F, 0x03, 0x59, 0x28, 0x75, 0x5D, 0x23, 0x28,
	0x11, 0x18, 0x5D, 0x15, 0x05, 0x5B, 0x30, 0x1C, 0x38, 0x1F, 0x1F, 0x07,
	0x19, 0x24, 0x05, 0x04, 0x06, 0x07, 0x57, 0x37, 0x3D, 0x0E, 0x07, 0x18,
	0x09, 0x09, 0x37, 0x21, 0x11, 0x37, 0x53, 0x31, 0x22, 0x13, 0x2B, 0x3D,
	0x2F, 0x15, 0x57, 0x08, 0x3D, 0x29, 0x29, 0x38, 0x0D, 0x33, 0x04, 0x3F,
	0x04, 0x2C, 0x0C, 0x3B, 0x29, 0x2C, 0x0C, 0x1D, 0x33, 0x29, 0x2E, 0x5C,
	0x03, 0x11, 0x00, 0x19, 0x34, 0x27, 0x27, 0x39, 0x14, 0x3F, 0x0D, 0x0B,
	0x5A, 0x2D, 0x58, 0x0C, 0x72, 0x58, 0x11, 0x2D, 0x2F, 0x2E, 0x1E, 0x29,
	0x59, 0x31, 0x20, 0x0D, 0x04, 0x0F, 0x1A, 0x33, 0x54, 0x4A, 0x1B, 0x40,
	0x0B, 0x54, 0x50, 0x20, 0x1D, 0x10, 0x2F, 0x0A, 0x59, 0x19, 0x21, 0x36,
	0x2B, 0x14, 0x1B, 0x08, 0x5F, 0x19, 0x3D, 0x05, 0x2F, 0x25, 0x17, 0x1F,
	0x3B, 0x76, 0x3A, 0x34, 0x38, 0x0E, 0x2B, 0x55, 0x39, 0x2D, 0x1A, 0x71,
	0x39, 0x0C, 0x45, 0x2C, 0x07, 0x23, 0x38, 0x39, 0x3C, 0x7B, 0x1C, 0x57,
	0x23, 0x21, 0x2E, 0x39, 0x06, 0x03, 0x39, 0x77, 0x5C, 0x15, 0x00, 0x0D,
	0x2E, 0x34, 0x30, 0x34, 0x53, 0x2C, 0x04, 0x51, 0x58, 0x03, 0x24, 0x5D,
	0x0B, 0x3B, 0x2D, 0x28, 0x5B, 0x0C, 0x3D, 0x00, 0x03, 0x34, 0x25, 0x05,
	0x04, 0x7B, 0x01, 0x12, 0x1F, 0x1A, 0x30, 0x43, 0x10, 0x05, 0x25, 0x38,
	0x2E, 0x22, 0x3C, 0x20, 0x0F, 0x58, 0x1B, 0x28, 0x3D, 0x31, 0x0B, 0x33,
	0x04, 0x5F, 0x03, 0x5F, 0x04, 0x07, 0x5D, 0x38, 0x3D, 0x2D, 0x36, 0x1E,
	0x0D, 0x1A, 0x56, 0x39, 0x25, 0x20, 0x00, 0x2D, 0x3B, 0x01, 0x2F, 0x3B,
	0x4A, 0x1C, 0x3A, 0x13, 0x01, 0x1B, 0x29, 0x02, 0x72, 0x03, 0x26, 0x0D,
	0x2E, 0x2F, 0x1C, 0x13, 0x07, 0x1B, 0x1A, 0x58, 0x08, 0x05, 0x31, 0x30,
	0x18, 0x02, 0x1F, 0x03, 0x34, 0x29, 0x13, 0x38, 0x19, 0x27, 0x5F, 0x0E,
	0x36, 0x52, 0x17, 0x3F, 0x50, 0x57, 0x02, 0x7A, 0x09, 0x23, 0x36, 0x44,
	0x36, 0x25, 0x39, 0x59, 0x3F, 0x27, 0x26, 0x2D, 0x18, 0x3D, 0x10, 0x1E,
	0x27, 0x1A, 0x19, 0x37, 0x05, 0x0D, 0x59, 0x38, 0x36, 0x34, 0x35, 0x39,
	0x40, 0x33, 0x05, 0x0F, 0x19, 0x3D, 0x34, 0x28, 0x36, 0x03, 0x31, 0x24,
	0x09, 0x54, 0x18, 0x28, 0x18, 0x02, 0x39, 0x3E, 0x38, 0x36, 0x0E, 0x06,
	0x5E, 0x18, 0x34, 0x03, 0x35, 0x2B, 0x0E, 0x7B, 0x1F, 0x2A, 0x38, 0x3C,
	0x35, 0x43, 0x33, 0x01, 0x38, 0x00, 0x0A, 0x24, 0x21, 0x01, 0x70, 0x0D,
	0x2A, 0x18, 0x28, 0x1B, 0x55, 0x32, 0x5A, 0x28, 0x36, 0x38, 0x2D, 0x2F,
	0x5F, 0x73, 0x36, 0x15, 0x02, 0x23, 0x09, 0x27, 0x54, 0x05, 0x24, 0x2B,
	0x36, 0x31, 0x37, 0x1C, 0x16, 0x55, 0x04, 0x1B, 0x18, 0x2C, 0x0E, 0x37,
	0x3B, 0x2C, 0x7B, 0x1B, 0x15, 0x03, 0x2C, 0x10, 0x01, 0x04, 0x3B, 0x18,
	0x08, 0x0D, 0x09, 0x23, 0x1E, 0x20, 0x2E, 0x36, 0x0C, 0x01, 0x21, 0x55,
	0x2A, 0x19, 0x0D, 0x11, 0x0D, 0x31, 0x3D, 0x29, 0x20, 0x09, 0x0D, 0x24,
	0x33, 0x7B, 0x36, 0x59, 0x5E, 0x22, 0x32, 0x5F, 0x09, 0x2C, 0x3A, 0x12,
	0x1C, 0x02, 0x2D, 0x38, 0x77, 0x24, 0x57, 0x0B, 0x32, 0x38, 0x20, 0x31,
	0x1F, 0x03, 0x69, 0x55, 0x27, 0x28, 0x22, 0x11, 0x2F, 0x37, 0x29, 0x39,
	0x32, 0x05, 0x32, 0x26, 0x04, 0x18, 0x59, 0x19, 0x41, 0x2D, 0x6D, 0x1A,
	0x12, 0x25, 0x5C, 0x26, 0x58, 0x17, 0x34, 0x3E, 0x21, 0x5D, 0x54, 0x29,
	0x08, 0x2C, 0x03, 0x36, 0x25, 0x22, 0x35, 0x1F, 0x26, 0x17, 0x03, 0x0C,
	0x5E, 0x02, 0x19, 0x5F, 0x1B, 0x3B, 0x32, 0x24, 0x0E, 0x73, 0x0D, 0x09,
	0x3A, 0x0A, 0x77, 0x34, 0x28, 0x57, 0x58, 0x76, 0x18, 0x0F, 0x16, 0x2A,
	0x2E, 0x3E, 0x2E, 0x16, 0x39, 0x26, 0x22, 0x33, 0x36, 0x33, 0x3B, 0x0B,
	0x51, 0x0F, 0x5D, 0x15, 0x21, 0x51, 0x17, 0x20, 0x07, 0x09, 0x19, 0x01,
	0x52, 0x1A, 0x1F, 0x32, 0x01, 0x3E, 0x74, 0x1D, 0x00, 0x02, 0x39, 0x17,
	0x14, 0x26, 0x0A, 0x0C, 0x1B, 0x14, 0x33, 0x18, 0x2F, 0x05, 0x1C, 0x33,
	0x5B, 0x5E, 0x11, 0x03, 0x54, 0x26, 0x12, 0x75, 0x07, 0x33, 0x08, 0x09,
	0x0F, 0x02, 0x2A, 0x08, 0x5B, 0x2F, 0x1D, 0x05, 0x17, 0x09, 0x0E, 0x2E,
	0x32, 0x2A, 0x5B, 0x2E, 0x23, 0x38, 0x2D, 0x27, 0x16, 0x25, 0x55, 0x05,
	0x2C, 0x11, 0x59, 0x13, 0x5C, 0x5F, 0x2A, 0x5B, 0x19, 0x1A, 0x32, 0x11,
	0x39, 0x50, 0x24, 0x2E, 0x23, 0x2F, 0x31, 0x06, 0x2A, 0x74, 0x18, 0x09,
	0x18, 0x31, 0x07, 0x38, 0x2F, 0x0F, 0x25, 0x11, 0x1D, 0x58, 0x25, 0x26,
	0x36, 0x3A, 0x26, 0x39, 0x19, 0x31, 0x09, 0x10, 0x41, 0x23, 0x11, 0x36,
	0x04, 0x3A, 0x3C, 0x35, 0x1E, 0x26, 0x59, 0x1A, 0x2D, 0x21, 0x0A, 0x0F,
	0x32, 0x31, 0x02, 0x58, 0x24, 0x44, 0x37, 0x2E, 0x3B, 0x04, 0x1D, 0x70,
	0x29, 0x05, 0x37, 0x1D, 0x77, 0x04, 0x32, 0x3C, 0x21, 0x13, 0x19, 0x35,
	0x5E, 0x53, 0x09, 0x06, 0x3B, 0x2A, 0x38, 0x05, 0x24, 0x02, 0x56, 0x02,
	0x29, 0x5E, 0x4E, 0x2D, 0x05, 0x77, 0x24, 0x05, 0x24, 0x25, 0x2F, 0x23,
	0x2A, 0x0D, 0x1C, 0x21, 0x3B, 0x36, 0x1B, 0x5A, 0x37, 0x28, 0x32, 0x36,
	0x5C, 0x09, 0x35, 0x51, 0x39, 0x5D, 0x16, 0x1C, 0x27, 0x05, 0x24, 0x2E,
	0x3F, 0x2B, 0x3B, 0x5F, 0x35, 0x05, 0x13, 0x23, 0x5C, 0x32, 0x03, 0x25,
	0x02, 0x58, 0x05, 0x3E, 0x4A, 0x0C, 0x52, 0x31, 0x29, 0x08, 0x0F, 0x5E,
	0x0C, 0x39, 0x0D, 0x5B, 0x1F, 0x2B, 0x3E, 0x28, 0x1C, 0x29, 0x1B, 0x03,
	0x50, 0x21, 0x0F, 0x08, 0x08, 0x13, 0x45, 0x09, 0x37, 0x16, 0x2A, 0x57,
	0x1D, 0x04, 0x5E, 0x23, 0x37, 0x03, 0x24, 0x01, 0x56, 0x08, 0x06, 0x27,
	0x3B, 0x0F, 0x25, 0x19, 0x76, 0x2D, 0x0B, 0x3E, 0x3F, 0x7B, 0x55, 0x2D,
	0x39, 0x1E, 0x32, 0x34, 0x2E, 0x29, 0x2C, 0x69, 0x15, 0x04, 0x22, 0x0A,
	0x20, 0x1F, 0x56, 0x2C, 0x2C, 0x28, 0x1C, 0x36, 0x59, 0x24, 0x20, 0x01,
	0x0B, 0x24, 0x11, 0x2A, 0x07, 0x23, 0x09, 0x1A, 0x2D, 0x22, 0x56, 0x0A,
	0x2C, 0x2B, 0x2D, 0x05, 0x23, 0x18, 0x23, 0x3F, 0x17, 0x2A, 0x52, 0x71,
	0x18, 0x09, 0x1D, 0x1B, 0x16, 0x1D, 0x24, 0x02, 0x5E, 0x0A, 0x5B, 0x17,
	0x2A, 0x19, 0x76, 0x47, 0x52, 0x58, 0x11, 0x13, 0x55, 0x13, 0x1F, 0x11,
	0x7B, 0x58, 0x38, 0x1F, 0x5D, 0x0F, 0x5C, 0x2D, 0x2B, 0x0E, 0x26, 0x14,
	0x58, 0x01, 0x2C, 0x16, 0x2B, 0x16, 0x2C, 0x19, 0x31, 0x06, 0x31, 0x02,
	0x5B, 0x14, 0x27, 0x0C, 0x1A, 0x11, 0x32, 0x02, 0x4A, 0x09, 0x5B, 0x15,
	0x0E, 0x2F, 0x39, 0x1B, 0x30, 0x2B, 0x2F, 0x0F, 0x01, 0x00, 0x18, 0x08,
	0x14, 0x04, 0x17, 0x5C, 0x06, 0x18, 0x5E, 0x17, 0x2F, 0x2C, 0x1D, 0x38,
	0x77, 0x02, 0x06, 0x2B, 0x33, 0x21, 0x1E, 0x22, 0x59, 0x05, 0x1A, 0x3D,
	0x04, 0x02, 0x38, 0x26, 0x36, 0x0D, 0x09, 0x1E, 0x2B, 0x2F, 0x06, 0x2A,
	0x19, 0x72, 0x2D, 0x12, 0x0D, 0x09, 0x26, 0x1D, 0x2B, 0x1D, 0x3D, 0x18,
	0x5D, 0x04, 0x01, 0x59, 0x38, 0x3E, 0x52, 0x0B, 0x40, 0x18, 0x06, 0x0F,
	0x0F, 0x3C, 0x08, 0x3F, 0x33, 0x45, 0x12, 0x35, 0x3C, 0x50, 0x5C, 0x52,
	0x04, 0x27, 0x14, 0x19, 0x05, 0x23, 0x1C, 0x55, 0x3F, 0x12, 0x1B, 0x19,
	0x09, 0x39, 0x3D, 0x25, 0x55, 0x37, 0x28, 0x25, 0x0A, 0x09, 0x05, 0x2F,
	0x08, 0x10, 0x3F, 0x27, 0x36, 0x0C, 0x2C, 0x04, 0x57, 0x0D, 0x1F, 0x0F,
	0x19, 0x17, 0x3B, 0x2C, 0x00, 0x1B, 0x34, 0x0D, 0x53, 0x70, 0x54, 0x35,
	0x04, 0x2C, 0x7A, 0x55, 0x23, 0x34, 0x3E, 0x74, 0x26, 0x2B, 0x34, 0x00,
	0x77, 0x55, 0x36, 0x00, 0x13, 0x11, 0x04, 0x02, 0x58, 0x11, 0x38, 0x14,
	0x10, 0x1D, 0x11, 0x2B, 0x2E, 0x54, 0x02, 0x3E, 0x24, 0x19, 0x29, 0x01,
	0x21, 0x05, 0x5F, 0x00, 0x25, 0x06, 0x0A, 0x19, 0x07, 0x00, 0x3A, 0x04,
	0x38, 0x25, 0x04, 0x3F, 0x7A, 0x35, 0x51, 0x5E, 0x5E, 0x17, 0x3B, 0x05,
	0x1A, 0x24, 0x11, 0x43, 0x29, 0x38, 0x25, 0x23, 0x23, 0x54, 0x5F, 0x2D,
	0x10, 0x38, 0x20, 0x5B, 0x33, 0x17, 0x14, 0x2B, 0x28, 0x58, 0x0F, 0x5A,
	0x11, 0x20, 0x01, 0x2D, 0x43, 0x36, 0x06, 0x1B, 0x2C, 0x07, 0x50, 0x3D,
	0x38, 0x18, 0x43, 0x1B, 0x29, 0x53, 0x35, 0x1C, 0x13, 0x0F, 0x04, 0x70,
	0x22, 0x0E, 0x19, 0x06, 0x32, 0x0E, 0x13, 0x1C, 0x03, 0x11, 0x25, 0x13,
	0x06, 0x3E, 0x28, 0x1A, 0x37, 0x20, 0x28, 0x23, 0x3C, 0x22, 0x05, 0x28,
	0x1B, 0x2D, 0x4E, 0x3A, 0x3E, 0x03, 0x43, 0x25, 0x39, 0x3F, 0x27, 0x35,
	0x20, 0x17, 0x21, 0x16, 0x1E, 0x14, 0x1C, 0x1E, 0x73, 0x0B, 0x02, 0x59,
	0x22, 0x17, 0x3B, 0x55, 0x41, 0x3D, 0x38, 0x35, 0x12, 0x36, 0x3D, 0x38,
	0x16, 0x0C, 0x5B, 0x38, 0x23, 0x55, 0x56, 0x0F, 0x28, 0x05, 0x1B, 0x0A,
	0x21, 0x3B, 0x23, 0x36, 0x0F, 0x1C, 0x12, 0x0F, 0x07, 0x14, 0x17, 0x1C,
	0x2C, 0x3F, 0x0D, 0x5F, 0x26, 0x0A, 0x34, 0x2C, 0x3F, 0x5A, 0x21, 0x29,
	0x54, 0x1A, 0x12, 0x34, 0x38, 0x14, 0x0B, 0x1E, 0x2B, 0x15, 0x39, 0x0B,
	0x25, 0x0C, 0x20, 0x11, 0x26, 0x1B, 0x37, 0x18, 0x16, 0x04, 0x19, 0x70,
	0x3B, 0x2F, 0x29, 0x04, 0x25, 0x15, 0x14, 0x1A, 0x0E, 0x30, 0x2A, 0x04,
	0x1D, 0x1E, 0x18, 0x22, 0x09, 0x28, 0x0A, 0x6D, 0x1C, 0x10, 0x28, 0x00,
	0x31, 0x3B, 0x4A, 0x1E, 0x3A, 0x3B, 0x3A, 0x37, 0x26, 0x3F, 0x37, 0x5C,
	0x24, 0x5C, 0x5D, 0x36, 0x02, 0x39, 0x3F, 0x2D, 0x2E, 0x36, 0x57, 0x3B,
	0x09, 0x09, 0x5F, 0x08, 0x02, 0x29, 0x0D, 0x5E, 0x26, 0x56, 0x53, 0x71,
	0x36, 0x00, 0x19, 0x1E, 0x03, 0x1C, 0x55, 0x1F, 0x13, 0x1A, 0x27, 0x2B,
	0x39, 0x12, 0x06, 0x34, 0x52, 0x14, 0x24, 0x10, 0x1E, 0x0F, 0x0F, 0x19,
	0x0B, 0x25, 0x30, 0x1B, 0x2E, 0x37, 0x02, 0x17, 0x58, 0x01, 0x13, 0x0E,
	0x2F, 0x3A, 0x22, 0x0D, 0x3A, 0x37, 0x3A, 0x07, 0x72, 0x55, 0x19, 0x09,
	0x1E, 0x77, 0x18, 0x26, 0x25, 0x3A, 0x7A, 0x43, 0x55, 0x58, 0x25, 0x13,
	0x18, 0x03, 0x5D, 0x05, 0x75, 0x15, 0x4E, 0x05, 0x26, 0x0B, 0x36, 0x54,
	0x37, 0x40, 0x74, 0x5B, 0x59, 0x37, 0x5D, 0x21, 0x38, 0x0B, 0x21, 0x1A,
	0x6D, 0x39, 0x08, 0x23, 0x3D, 0x73, 0x29, 0x4A, 0x1D, 0x26, 0x15, 0x03,
	0x05, 0x0D, 0x5B, 0x29, 0x20, 0x56, 0x22, 0x1B, 0x73, 0x2B, 0x2C, 0x1C,
	0x29, 0x21, 0x3B, 0x22, 0x17, 0x07, 0x27, 0x07, 0x27, 0x16, 0x0A, 0x10,
	0x39, 0x10, 0x36, 0x27, 0x20, 0x5A, 0x06, 0x5F, 0x59, 0x13, 0x0A, 0x53,
	0x25, 0x03, 0x2A, 0x5D, 0x1B, 0x03, 0x05, 0x0E, 0x27, 0x12, 0x36, 0x1E,
	0x15, 0x06, 0x03, 0x1B, 0x21, 0x2C, 0x08, 0x13, 0x2B, 0x25, 0x2A, 0x0D,
	0x57, 0x0F, 0x39, 0x30, 0x3A, 0x29, 0x34, 0x25, 0x10, 0x5A, 0x31, 0x08,
	0x0D, 0x2A, 0x15, 0x1B, 0x2D, 0x2C, 0x0F, 0x15, 0x38, 0x3E, 0x58, 0x16,
	0x1E, 0x07, 0x1C, 0x25, 0x29, 0x0D, 0x38, 0x1F, 0x5C, 0x38, 0x2A, 0x05,
	0x0A, 0x0F, 0x24, 0x1C, 0x28, 0x0B, 0x1B, 0x17, 0x3E, 0x31, 0x18, 0x0E,
	0x18, 0x35, 0x3B, 0x29, 0x03, 0x32, 0x3C, 0x0A, 0x1E, 0x1E, 0x18, 0x5C,
	0x12, 0x2A, 0x01, 0x31, 0x34, 0x06, 0x0B, 0x5C, 0x14, 0x5A, 0x2E, 0x41,
	0x1C, 0x72, 0x58, 0x03, 0x41, 0x39, 0x04, 0x29, 0x0F, 0x39, 0x13, 0x10,
	0x2F, 0x36, 0x57, 0x27, 0x35, 0x3A, 0x53, 0x0A, 0x3C, 0x27, 0x27, 0x07,
	0x2F, 0x02, 0x76, 0x01, 0x16, 0x24, 0x27, 0x30, 0x16, 0x38, 0x5B, 0x32,
	0x05, 0x08, 0x22, 0x16, 0x06, 0x0A, 0x06, 0x26, 0x5B, 0x1A, 0x3A, 0x02,
	0x05, 0x37, 0x28, 0x2C, 0x09, 0x16, 0x0F, 0x22, 0x0D, 0x07, 0x11, 0x0D,
	0x07, 0x23, 0x0A, 0x0D, 0x59, 0x1E, 0x03, 0x19, 0x54, 0x1C, 0x0C, 0x28,
	0x14, 0x50, 0x3D, 0x12, 0x0F, 0x3E, 0x15, 0x22, 0x52, 0x0F, 0x20, 0x23,
	0x3D, 0x23, 0x36, 0x08, 0x50, 0x24, 0x1D, 0x34, 0x00, 0x31, 0x22, 0x3E,
	0x12, 0x3B, 0x2D, 0x09, 0x39, 0x33, 0x18, 0x05, 0x20, 0x2A, 0x20, 0x08,
	0x2B, 0x2B, 0x38, 0x7B, 0x5A, 0x34, 0x1A, 0x23, 0x76, 0x1D, 0x2B, 0x37,
	0x0F, 0x10, 0x18, 0x1B, 0x3E, 0x04, 0x26, 0x38, 0x14, 0x20, 0x06, 0x36,
	0x21, 0x4A, 0x1D, 0x3E, 0x1A, 0x55, 0x37, 0x16, 0x1E, 0x2A, 0x29, 0x0C,
	0x5B, 0x06, 0x13, 0x38, 0x30, 0x02, 0x27, 0x01, 0x01, 0x3B, 0x0D, 0x31,
	0x31, 0x5C, 0x4A, 0x3E, 0x08, 0x73, 0x5C, 0x2C, 0x5B, 0x5A, 0x28, 0x0D,
	0x0A, 0x37, 0x5D, 0x71, 0x08, 0x26, 0x5A, 0x19, 0x36, 0x29, 0x02, 0x1A,
	0x3D, 0x26, 0x14, 0x3B, 0x17, 0x01, 0x2A, 0x2A, 0x39, 0x03, 0x05, 0x00,
	0x22, 0x2A, 0x1A, 0x21, 0x04, 0x04, 0x4A, 0x09, 0x0E, 0x70, 0x09, 0x2D,
	0x22, 0x07, 0x29, 0x18, 0x26, 0x28, 0x29, 0x2C, 0x3D, 0x15, 0x1E, 0x11,
	0x0E, 0x08, 0x2A, 0x2F, 0x07, 0x7B, 0x5E, 0x17, 0x2A, 0x21, 0x0D, 0x04,
	0x18, 0x0B, 0x19, 0x72, 0x3C, 0x2B, 0x5B, 0x31, 0x29, 0x23, 0x0C, 0x36,
	0x2C, 0x0D, 0x03, 0x05, 0x16, 0x1A, 0x06, 0x3F, 0x24, 0x1B, 0x3C, 0x2E,
	0x3A, 0x14, 0x03, 0x26, 0x14, 0x07, 0x58, 0x5D, 0x13, 0x00, 0x5C, 0x37,
	0x39, 0x0A, 0x0D, 0x3E, 0x1B, 0x45, 0x03, 0x08, 0x3C, 0x50, 0x1E, 0x02,
	0x70, 0x1D, 0x13, 0x57, 0x33, 0x15, 0x59, 0x19, 0x3B, 0x19, 0x33, 0x36,
	0x51, 0x23, 0x38, 0x26, 0x3A, 0x38, 0x25, 0x26, 0x17, 0x1C, 0x04, 0x2A,
	0x39, 0x20, 0x43, 0x0A, 0x0B, 0x18, 0x21, 0x5C, 0x56, 0x25, 0x39, 0x74,
	0x55, 0x24, 0x24, 0x5C, 0x74, 0x00, 0x32, 0x0F, 0x1D, 0x74, 0x1D, 0x2C,
	0x59, 0x5D, 0x38, 0x05, 0x00, 0x21, 0x06, 0x3B, 0x1A, 0x37, 0x59, 0x40,
	0x0B, 0x3B, 0x53, 0x09, 0x26, 0x69, 0x59, 0x22, 0x5B, 0x59, 0x10, 0x39,
	0x0D, 0x3C, 0x1F, 0x14, 0x3F, 0x00, 0x1C, 0x25, 0x2F, 0x54, 0x2A, 0x5B,
	0x32, 0x2F, 0x14, 0x0F, 0x0C, 0x20, 0x26, 0x14, 0x05, 0x18, 0x38, 0x15,
	0x5B, 0x2E, 0x59, 0x09, 0x77, 0x2D, 0x23, 0x04, 0x25, 0x2E, 0x2A, 0x54,
	0x1C, 0x3E, 0x21, 0x19, 0x33, 0x3C, 0x1A, 0x14, 0x1E, 0x50, 0x14, 0x13,
	0x38, 0x07, 0x02, 0x39, 0x1B, 0x3A, 0x1A, 0x35, 0x0A, 0x0E, 0x07, 0x01,
	0x04, 0x5B, 0x08, 0x2F, 0x00, 0x22, 0x5B, 0x5C, 0x05, 0x16, 0x14, 0x2B,
	0x18, 0x2A, 0x36, 0x32, 0x3E, 0x0A, 0x72, 0x54, 0x19, 0x09, 0x26, 0x13,
	0x08, 0x19, 0x14, 0x21, 0x71, 0x35, 0x50, 0x14, 0x00, 0x2A, 0x25, 0x57,
	0x0C, 0x1A, 0x33, 0x0B, 0x14, 0x56, 0x2E, 0x28, 0x1F, 0x51, 0x3D, 0x1A,
	0x15, 0x47, 0x23, 0x27, 0x0E, 0x16, 0x5B, 0x11, 0x5F, 0x04, 0x1A, 0x07,
	0x37, 0x2C, 0x09, 0x6D, 0x22, 0x23, 0x29, 0x0E, 0x04, 0x16, 0x2F, 0x29,
	0x05, 0x0A, 0x5E, 0x07, 0x17, 0x09, 0x2C, 0x3E, 0x28, 0x04, 0x26, 0x2E,
	0x38, 0x39, 0x14, 0x3B, 0x7A, 0x20, 0x39, 0x0A, 0x53, 0x25, 0x21, 0x05,
	0x2D, 0x58, 0x69, 0x3C, 0x34, 0x23, 0x07, 0x01, 0x5D, 0x34, 0x17, 0x3E,
	0x7B, 0x38, 0x08, 0x3D, 0x19, 0x24, 0x1C, 0x0A, 0x1F, 0x1D, 0x2C, 0x36,
	0x28, 0x0D, 0x5F, 0x00, 0x23, 0x2D, 0x19, 0x13, 0x12, 0x55, 0x53, 0x24,
	0x19, 0x0D, 0x1E, 0x4A, 0x5C, 0x1D, 0x38, 0x5F, 0x04, 0x1D, 0x24, 0x73,
	0x3A, 0x30, 0x0F, 0x2C, 0x27, 0x23, 0x0C, 0x41, 0x39, 0x16, 0x21, 0x2C,
	0x5C, 0x5C, 0x11, 0x3D, 0x27, 0x24, 0x06, 0x1B, 0x39, 0x56, 0x0C, 0x08,
	0x36, 0x43, 0x56, 0x0A, 0x3F, 0x3A, 0x28, 0x53, 0x36, 0x5D, 0x12, 0x0D,
	0x32, 0x1A, 0x31, 0x0D, 0x5C, 0x08, 0x3E, 0x52, 0x00, 0x34, 0x27, 0x3A,
	0x0C, 0x3B, 0x2F, 0x13, 0x24, 0x1B, 0x2B, 0x5F, 0x11, 0x24, 0x03, 0x70,
	0x43, 0x30, 0x59, 0x07, 0x06, 0x35, 0x30, 0x06, 0x18, 0x2D, 0x3A, 0x07,
	0x07, 0x5A, 0x0C, 0x0F, 0x15, 0x26, 0x24, 0x32, 0x58, 0x10, 0x2A, 0x3D,
	0x75, 0x29, 0x50, 0x17, 0x11, 0x7B, 0x06, 0x14, 0x3B, 0x0E, 0x31, 0x5A,
	0x26, 0x0B, 0x0D, 0x09, 0x06, 0x13, 0x24, 0x44, 0x0B, 0x5C, 0x53, 0x22,
	0x5B, 0x37, 0x19, 0x0D, 0x1F, 0x39, 0x12, 0x07, 0x50, 0x3B, 0x27, 0x2C,
	0x39, 0x0E, 0x21, 0x5A, 0x36, 0x22, 0x11, 0x0C, 0x3A, 0x7B, 0x09, 0x34,
	0x20, 0x2A, 0x2E, 0x1E, 0x0F, 0x04, 0x40, 0x20, 0x14, 0x22, 0x23, 0x5C,
	0x00, 0x0F, 0x32, 0x0D, 0x59, 0x25, 0x2B, 0x55, 0x3A, 0x3F, 0x0C, 0x3B,
	0x26, 0x3F, 0x01, 0x18, 0x59, 0x56, 0x3A, 0x22, 0x75, 0x3F, 0x03, 0x5F,
	0x32, 0x15, 0x3C, 0x2C, 0x21, 0x26, 0x27, 0x1A, 0x53, 0x1B, 0x02, 0x0E,
	0x3A, 0x55, 0x3D, 0x0D, 0x0E, 0x3A, 0x32, 0x0D, 0x39, 0x75, 0x3E, 0x08,
	0x1F, 0x08, 0x3B, 0x0F, 0x28, 0x57, 0x32, 0x20, 0x21, 0x58, 0x25, 0x5E,
	0x0D, 0x1D, 0x14, 0x03, 0x1B, 0x0E, 0x5A, 0x36, 0x29, 0x5A, 0x7A, 0x00,
	0x19, 0x58, 0x31, 0x10, 0x59, 0x04, 0x1C, 0x00, 0x33, 0x1C, 0x18, 0x3F,
	0x24, 0x36, 0x34, 0x00, 0x58, 0x20, 0x20, 0x25, 0x23, 0x29, 0x32, 0x05,
	0x1A, 0x35, 0x22, 0x04, 0x75, 0x2B, 0x03, 0x0C, 0x5B, 0x72, 0x34, 0x35,
	0x2F, 0x20, 0x03, 0x55, 0x32, 0x0A, 0x1A, 0x21, 0x1A, 0x59, 0x07, 0x1B,
	0x13, 0x43, 0x0E, 0x58, 0x12, 0x10, 0x58, 0x4A, 0x1C, 0x13, 0x11, 0x5A,
	0x10, 0x1E, 0x08, 0x28, 0x18, 0x06, 0x59, 0x1B, 0x3B, 0x5E, 0x08, 0x2B,
	0x24, 0x29, 0x1E, 0x2B, 0x1C, 0x1D, 0x30, 0x5B, 0x2B, 0x17, 0x01, 0x15,
	0x0E, 0x2E, 0x28, 0x18, 0x34, 0x3F, 0x15, 0x5D, 0x38, 0x14, 0x1C, 0x15,
	0x5D, 0x32, 0x37, 0x35, 0x4A, 0x08, 0x3D, 0x2A, 0x36, 0x32, 0x5B, 0x19,
	0x1A, 0x0D, 0x55, 0x5D, 0x0F, 0x06, 0x03, 0x22, 0x25, 0x02, 0x0F, 0x35,
	0x13, 0x3B, 0x04, 0x06, 0x02, 0x15, 0x08, 0x5D, 0x28, 0x2A, 0x2C, 0x16,
	0x3D, 0x1B, 0x09, 0x55, 0x45, 0x24, 0x0F, 0x00, 0x53, 0x59, 0x0E, 0x73,
	0x5F, 0x05, 0x1C, 0x31, 0x6D, 0x18, 0x2F, 0x18, 0x3F, 0x00, 0x39, 0x08,
	0x07, 0x0D, 0x2E, 0x55, 0x2A, 0x5F, 0x0E, 0x37, 0x39, 0x30, 0x1A, 0x23,
	0x72, 0x01, 0x2F, 0x25, 0x09, 0x71, 0x04, 0x29, 0x01, 0x02, 0x16, 0x0E,
	0x0F, 0x24, 0x22, 0x07, 0x1F, 0x33, 0x29, 0x58, 0x71, 0x43, 0x19, 0x41,
	0x09, 0x23, 0x26, 0x27, 0x17, 0x1C, 0x7F, 0x51]

	data = xorcrypt(data)
	data = base64.decode(data.bytestr())
	data = zlib.decompress(data)!

	return data
}

pub fn getdata() []u8 {
	return decompress() or {
		println('Error')
		exit(1)
	}
}